--//////////////////////////////////////////////////////////////////////////////
-- Project Name:	CoCo3FPGA Version 4.0
-- File Name:		coco_rom.vhd
--
-- CoCo3 in an FPGA
--
-- Revision: 4.0 07/10/16
--//////////////////////////////////////////////////////////////////////////////
--
-- CPU section copyrighted by John Kent
-- The FDC co-processor copyrighted Daniel Wallner.
-- SDRAM Controller copyrighted by XESS Corp.
--
--//////////////////////////////////////////////////////////////////////////////
--
-- Color Computer 3 compatible system on a chip
--
-- Version : 4.1.2
--
-- Copyright (c) 2008 Gary Becker (gary_l_becker@yahoo.com)
--
-- All rights reserved
--
-- Redistribution and use in source and synthezised forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- Redistributions of source code must retain the above copyright notice,
-- this list of conditions and the following disclaimer.
--																		   
-- Redistributions in synthesized form must reproduce the above copyright
-- notice, this list of conditions and the following disclaimer in the
-- documentation and/or other materials provided with the distribution.
--
-- Neither the name of the author nor the names of other contributors may
-- be used to endorse or promote products derived from this software without
-- specific prior written permission.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
--
-- Please report bugs to the author, but before you do so, please
-- make sure that this is not a derivative work and that
-- you have the latest version of this file.
--
-- The latest version of this file can be found at:
--      http://groups.yahoo.com/group/CoCo3FPGA
--
-- File history :
--
--  1.0			Full Release
--  2.0			Partial Release
--  3.0			Full Release
--  3.0.0.1		Update to fix DoD interrupt issue
--	3.0.1.0		Update to fix 32/40 CoCO3 Text issue and add 2 Meg max memory
--	4.0.X.X		Full Release
--	4.1.2.X		Fixed 6502 code for drivewire, removed timer, fixed 6551 baud 
--				rate (& DE2-115 compiler symbol)
--//////////////////////////////////////////////////////////////////////////////
-- Gary Becker
-- gary_L_becker@yahoo.com
--//////////////////////////////////////////////////////////////////////////////
--//////////////////////////////////////////////////////////////////////////////
-- DE2-115 Conversion by Stan Hodge
-- shodgefamily@yahoo.com
--//////////////////////////////////////////////////////////////////////////////
-- MISTer conversion work by Stan Hodge and Alan Steremberg

-- generated with romgen v3.0 by MikeJ

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity COCO_ROM is
  port (
    ADDR        : in    std_logic_vector(15 downto 0);
    DATA        : out   std_logic_vector(7 downto 0);
	 CLK : in std_logic;
	 WR_ADDR : in std_logic_vector(15 downto 0);
	 WR_DATA : in std_logic_vector(7 downto 0);
	 WR : in std_logic
    );
end;

architecture RTL of COCO_ROM is


  type ROM_ARRAY is array(0 to 65535) of std_logic_vector(7 downto 0);
  signal ROM : ROM_ARRAY := (
    x"45",x"58",x"8E",x"80",x"DE",x"CE",x"01",x"2A", -- 0x0000
    x"C6",x"0A",x"BD",x"A5",x"9A",x"8E",x"B2",x"77", -- 0x0008
    x"AF",x"43",x"AF",x"48",x"8E",x"89",x"4C",x"BF", -- 0x0010
    x"01",x"0D",x"9E",x"8A",x"BF",x"01",x"12",x"BD", -- 0x0018
    x"82",x"9C",x"CC",x"2C",x"05",x"DD",x"E6",x"8E", -- 0x0020
    x"01",x"3E",x"9F",x"B0",x"CE",x"B4",x"4A",x"C6", -- 0x0028
    x"0A",x"EF",x"81",x"5A",x"26",x"FB",x"86",x"7E", -- 0x0030
    x"B7",x"01",x"9A",x"8E",x"82",x"B9",x"BF",x"01", -- 0x0038
    x"9B",x"B7",x"01",x"8B",x"8E",x"88",x"46",x"BF", -- 0x0040
    x"01",x"8C",x"B7",x"01",x"97",x"8E",x"87",x"E5", -- 0x0048
    x"BF",x"01",x"98",x"B7",x"01",x"79",x"8E",x"8E", -- 0x0050
    x"90",x"BF",x"01",x"7A",x"B7",x"01",x"91",x"8E", -- 0x0058
    x"88",x"F0",x"BF",x"01",x"92",x"B7",x"01",x"6A", -- 0x0060
    x"8E",x"8C",x"F1",x"BF",x"01",x"6B",x"B7",x"01", -- 0x0068
    x"67",x"8E",x"82",x"73",x"BF",x"01",x"68",x"B7", -- 0x0070
    x"01",x"76",x"8E",x"82",x"86",x"BF",x"01",x"77", -- 0x0078
    x"B7",x"01",x"A3",x"8E",x"83",x"04",x"BF",x"01", -- 0x0080
    x"A4",x"B7",x"01",x"94",x"8E",x"82",x"9C",x"BF", -- 0x0088
    x"01",x"95",x"B7",x"01",x"1D",x"8E",x"84",x"89", -- 0x0090
    x"BF",x"01",x"1E",x"BD",x"96",x"E6",x"B6",x"FF", -- 0x0098
    x"03",x"8A",x"01",x"B7",x"FF",x"03",x"8E",x"44", -- 0x00A0
    x"4B",x"BC",x"C0",x"00",x"10",x"27",x"3F",x"52", -- 0x00A8
    x"1C",x"AF",x"8E",x"80",x"E7",x"BD",x"B9",x"9C", -- 0x00B0
    x"8E",x"80",x"C0",x"9F",x"72",x"7E",x"A0",x"E2", -- 0x00B8
    x"FF",x"0F",x"E3",x"0F",x"E4",x"B6",x"FF",x"03", -- 0x00C0
    x"8A",x"01",x"B7",x"FF",x"03",x"7E",x"A0",x"E8", -- 0x00C8
    x"96",x"68",x"4C",x"27",x"08",x"1F",x"20",x"93", -- 0x00D0
    x"19",x"D3",x"A6",x"DD",x"A6",x"39",x"19",x"81", -- 0x00D8
    x"83",x"81",x"3C",x"0E",x"82",x"1E",x"81",x"68", -- 0x00E0
    x"45",x"58",x"54",x"45",x"4E",x"44",x"45",x"44", -- 0x00E8
    x"20",x"43",x"4F",x"4C",x"4F",x"52",x"20",x"42", -- 0x00F0
    x"41",x"53",x"49",x"43",x"20",x"32",x"2E",x"30", -- 0x00F8
    x"0D",x"43",x"4F",x"50",x"52",x"2E",x"20",x"31", -- 0x0100
    x"39",x"38",x"32",x"2C",x"20",x"31",x"39",x"38", -- 0x0108
    x"36",x"20",x"42",x"59",x"20",x"54",x"41",x"4E", -- 0x0110
    x"44",x"59",x"20",x"20",x"0D",x"55",x"4E",x"44", -- 0x0118
    x"45",x"52",x"20",x"4C",x"49",x"43",x"45",x"4E", -- 0x0120
    x"53",x"45",x"20",x"46",x"52",x"4F",x"4D",x"20", -- 0x0128
    x"4D",x"49",x"43",x"52",x"4F",x"53",x"4F",x"46", -- 0x0130
    x"54",x"0D",x"0D",x"00",x"81",x"CB",x"22",x"08", -- 0x0138
    x"8E",x"81",x"F0",x"80",x"B5",x"7E",x"AD",x"D4", -- 0x0140
    x"81",x"FF",x"27",x"08",x"81",x"CD",x"23",x"15", -- 0x0148
    x"6E",x"9F",x"01",x"37",x"9D",x"9F",x"81",x"90", -- 0x0150
    x"10",x"27",x"05",x"7A",x"81",x"9F",x"10",x"27", -- 0x0158
    x"07",x"FE",x"BD",x"01",x"A0",x"7E",x"B2",x"77", -- 0x0160
    x"C1",x"42",x"23",x"04",x"6E",x"9F",x"01",x"3C", -- 0x0168
    x"C0",x"28",x"C1",x"10",x"22",x"07",x"34",x"04", -- 0x0170
    x"BD",x"B2",x"62",x"35",x"04",x"8E",x"82",x"57", -- 0x0178
    x"7E",x"B2",x"CE",x"44",x"45",x"CC",x"45",x"44", -- 0x0180
    x"49",x"D4",x"54",x"52",x"4F",x"CE",x"54",x"52", -- 0x0188
    x"4F",x"46",x"C6",x"44",x"45",x"C6",x"4C",x"45", -- 0x0190
    x"D4",x"4C",x"49",x"4E",x"C5",x"50",x"43",x"4C", -- 0x0198
    x"D3",x"50",x"53",x"45",x"D4",x"50",x"52",x"45", -- 0x01A0
    x"53",x"45",x"D4",x"53",x"43",x"52",x"45",x"45", -- 0x01A8
    x"CE",x"50",x"43",x"4C",x"45",x"41",x"D2",x"43", -- 0x01B0
    x"4F",x"4C",x"4F",x"D2",x"43",x"49",x"52",x"43", -- 0x01B8
    x"4C",x"C5",x"50",x"41",x"49",x"4E",x"D4",x"47", -- 0x01C0
    x"45",x"D4",x"50",x"55",x"D4",x"44",x"52",x"41", -- 0x01C8
    x"D7",x"50",x"43",x"4F",x"50",x"D9",x"50",x"4D", -- 0x01D0
    x"4F",x"44",x"C5",x"50",x"4C",x"41",x"D9",x"44", -- 0x01D8
    x"4C",x"4F",x"41",x"C4",x"52",x"45",x"4E",x"55", -- 0x01E0
    x"CD",x"46",x"CE",x"55",x"53",x"49",x"4E",x"C7", -- 0x01E8
    x"89",x"70",x"85",x"33",x"86",x"A7",x"86",x"A8", -- 0x01F0
    x"88",x"71",x"AF",x"89",x"93",x"BB",x"95",x"32", -- 0x01F8
    x"93",x"61",x"93",x"65",x"96",x"70",x"96",x"8B", -- 0x0200
    x"95",x"46",x"9E",x"9D",x"98",x"EC",x"97",x"55", -- 0x0208
    x"97",x"58",x"9C",x"B6",x"97",x"23",x"96",x"21", -- 0x0210
    x"9A",x"22",x"8C",x"18",x"8A",x"09",x"41",x"54", -- 0x0218
    x"CE",x"43",x"4F",x"D3",x"54",x"41",x"CE",x"45", -- 0x0220
    x"58",x"D0",x"46",x"49",x"D8",x"4C",x"4F",x"C7", -- 0x0228
    x"50",x"4F",x"D3",x"53",x"51",x"D2",x"48",x"45", -- 0x0230
    x"58",x"A4",x"56",x"41",x"52",x"50",x"54",x"D2", -- 0x0238
    x"49",x"4E",x"53",x"54",x"D2",x"54",x"49",x"4D", -- 0x0240
    x"45",x"D2",x"50",x"50",x"4F",x"49",x"4E",x"D4", -- 0x0248
    x"53",x"54",x"52",x"49",x"4E",x"47",x"A4",x"83", -- 0x0250
    x"B0",x"83",x"78",x"83",x"81",x"84",x"F2",x"85", -- 0x0258
    x"24",x"84",x"46",x"86",x"AC",x"84",x"80",x"8B", -- 0x0260
    x"DD",x"86",x"BE",x"87",x"7E",x"89",x"68",x"93", -- 0x0268
    x"39",x"87",x"4E",x"0D",x"6F",x"10",x"27",x"13", -- 0x0270
    x"33",x"34",x"04",x"D6",x"6F",x"C1",x"FD",x"35", -- 0x0278
    x"04",x"26",x"02",x"32",x"62",x"39",x"96",x"6F", -- 0x0280
    x"4C",x"26",x"FA",x"96",x"78",x"81",x"02",x"26", -- 0x0288
    x"F4",x"96",x"79",x"26",x"F0",x"0F",x"6F",x"32", -- 0x0290
    x"62",x"7E",x"A4",x"44",x"CC",x"BA",x"42",x"DD", -- 0x0298
    x"DF",x"86",x"02",x"97",x"E2",x"97",x"DE",x"48", -- 0x02A0
    x"97",x"E1",x"0F",x"E5",x"DC",x"8A",x"DD",x"E8", -- 0x02A8
    x"C6",x"80",x"DD",x"C7",x"C6",x"60",x"DD",x"C9", -- 0x02B0
    x"39",x"32",x"62",x"1C",x"AF",x"BD",x"AD",x"EB", -- 0x02B8
    x"9E",x"A6",x"9F",x"2F",x"A6",x"80",x"27",x"07", -- 0x02C0
    x"81",x"3A",x"27",x"25",x"7E",x"B2",x"77",x"A6", -- 0x02C8
    x"81",x"97",x"00",x"26",x"03",x"7E",x"AE",x"15", -- 0x02D0
    x"EC",x"80",x"DD",x"68",x"9F",x"A6",x"96",x"AF", -- 0x02D8
    x"27",x"0F",x"86",x"5B",x"BD",x"A2",x"82",x"96", -- 0x02E0
    x"68",x"BD",x"BD",x"CC",x"86",x"5D",x"BD",x"A2", -- 0x02E8
    x"82",x"9D",x"9F",x"1F",x"A9",x"81",x"98",x"27", -- 0x02F0
    x"1D",x"81",x"97",x"27",x"14",x"1F",x"9A",x"BD", -- 0x02F8
    x"AD",x"C6",x"20",x"B7",x"AE",x"62",x"8C",x"AC", -- 0x0300
    x"9D",x"26",x"05",x"8E",x"82",x"F1",x"AF",x"62", -- 0x0308
    x"39",x"BD",x"8C",x"62",x"20",x"A5",x"8D",x"02", -- 0x0310
    x"20",x"A1",x"9D",x"9F",x"81",x"4D",x"10",x"26", -- 0x0318
    x"21",x"2A",x"9D",x"9F",x"BD",x"A5",x"78",x"8D", -- 0x0320
    x"43",x"BF",x"01",x"E7",x"8D",x"3E",x"AC",x"62", -- 0x0328
    x"10",x"25",x"31",x"16",x"8D",x"36",x"BF",x"01", -- 0x0330
    x"E5",x"9D",x"A5",x"26",x"D3",x"86",x"02",x"9E", -- 0x0338
    x"8A",x"BD",x"A6",x"5F",x"0F",x"78",x"0C",x"7C", -- 0x0340
    x"BD",x"A7",x"D8",x"AE",x"64",x"9F",x"7E",x"86", -- 0x0348
    x"FF",x"97",x"7D",x"EC",x"62",x"93",x"7E",x"24", -- 0x0350
    x"05",x"32",x"66",x"7E",x"A4",x"91",x"10",x"83", -- 0x0358
    x"00",x"FF",x"24",x"03",x"5C",x"D7",x"7D",x"BD", -- 0x0360
    x"A7",x"F4",x"20",x"E1",x"BD",x"B2",x"6D",x"BD", -- 0x0368
    x"B7",x"3D",x"EE",x"E4",x"AF",x"E4",x"1F",x"35", -- 0x0370
    x"8E",x"83",x"AB",x"BD",x"B9",x"C2",x"7E",x"BF", -- 0x0378
    x"78",x"BD",x"BC",x"2F",x"0F",x"0A",x"8D",x"F6", -- 0x0380
    x"8E",x"00",x"4A",x"BD",x"BC",x"35",x"8E",x"00", -- 0x0388
    x"40",x"BD",x"BC",x"14",x"0F",x"54",x"96",x"0A", -- 0x0390
    x"8D",x"0C",x"0D",x"4F",x"10",x"27",x"36",x"F2", -- 0x0398
    x"8E",x"00",x"4A",x"7E",x"BB",x"8F",x"34",x"02", -- 0x03A0
    x"7E",x"BF",x"A6",x"81",x"49",x"0F",x"DA",x"A2", -- 0x03A8
    x"96",x"54",x"34",x"02",x"2A",x"02",x"8D",x"24", -- 0x03B0
    x"96",x"4F",x"34",x"02",x"81",x"81",x"25",x"05", -- 0x03B8
    x"8E",x"BA",x"C5",x"8D",x"DE",x"8E",x"83",x"E0", -- 0x03C0
    x"BD",x"BE",x"F0",x"35",x"02",x"81",x"81",x"25", -- 0x03C8
    x"06",x"8E",x"83",x"AB",x"BD",x"B9",x"B9",x"35", -- 0x03D0
    x"02",x"4D",x"2A",x"03",x"7E",x"BE",x"E9",x"39", -- 0x03D8
    x"0B",x"76",x"B3",x"83",x"BD",x"D3",x"79",x"1E", -- 0x03E0
    x"F4",x"A6",x"F5",x"7B",x"83",x"FC",x"B0",x"10", -- 0x03E8
    x"7C",x"0C",x"1F",x"67",x"CA",x"7C",x"DE",x"53", -- 0x03F0
    x"CB",x"C1",x"7D",x"14",x"64",x"70",x"4C",x"7D", -- 0x03F8
    x"B7",x"EA",x"51",x"7A",x"7D",x"63",x"30",x"88", -- 0x0400
    x"7E",x"7E",x"92",x"44",x"99",x"3A",x"7E",x"4C", -- 0x0408
    x"CC",x"91",x"C7",x"7F",x"AA",x"AA",x"AA",x"13", -- 0x0410
    x"81",x"00",x"00",x"00",x"00",x"03",x"7F",x"5E", -- 0x0418
    x"56",x"CB",x"79",x"80",x"13",x"9B",x"0B",x"64", -- 0x0420
    x"80",x"76",x"38",x"93",x"16",x"82",x"38",x"AA", -- 0x0428
    x"3B",x"20",x"80",x"35",x"04",x"F3",x"34",x"81", -- 0x0430
    x"35",x"04",x"F3",x"34",x"80",x"80",x"00",x"00", -- 0x0438
    x"00",x"80",x"31",x"72",x"17",x"F8",x"BD",x"BC", -- 0x0440
    x"6D",x"10",x"2F",x"2F",x"FD",x"8E",x"84",x"32", -- 0x0448
    x"96",x"4F",x"80",x"80",x"34",x"02",x"86",x"80", -- 0x0450
    x"97",x"4F",x"BD",x"B9",x"C2",x"8E",x"84",x"37", -- 0x0458
    x"BD",x"BB",x"8F",x"8E",x"BA",x"C5",x"BD",x"B9", -- 0x0460
    x"B9",x"8E",x"84",x"1D",x"BD",x"BE",x"F0",x"8E", -- 0x0468
    x"84",x"3C",x"BD",x"B9",x"C2",x"35",x"04",x"BD", -- 0x0470
    x"BD",x"99",x"8E",x"84",x"41",x"7E",x"BA",x"CA", -- 0x0478
    x"BD",x"BC",x"5F",x"8E",x"BE",x"C0",x"BD",x"BC", -- 0x0480
    x"14",x"27",x"67",x"4D",x"26",x"03",x"7E",x"BA", -- 0x0488
    x"3A",x"8E",x"00",x"4A",x"BD",x"BC",x"35",x"5F", -- 0x0490
    x"96",x"61",x"2A",x"10",x"BD",x"BC",x"EE",x"8E", -- 0x0498
    x"00",x"4A",x"96",x"61",x"BD",x"BC",x"A0",x"26", -- 0x04A0
    x"03",x"43",x"D6",x"01",x"BD",x"BC",x"4C",x"34", -- 0x04A8
    x"04",x"BD",x"84",x"46",x"8E",x"00",x"4A",x"BD", -- 0x04B0
    x"BA",x"CA",x"8D",x"36",x"35",x"02",x"46",x"10", -- 0x04B8
    x"25",x"3A",x"26",x"39",x"81",x"38",x"AA",x"3B", -- 0x04C0
    x"29",x"07",x"71",x"34",x"58",x"3E",x"56",x"74", -- 0x04C8
    x"16",x"7E",x"B3",x"1B",x"77",x"2F",x"EE",x"E3", -- 0x04D0
    x"85",x"7A",x"1D",x"84",x"1C",x"2A",x"7C",x"63", -- 0x04D8
    x"59",x"58",x"0A",x"7E",x"75",x"FD",x"E7",x"C6", -- 0x04E0
    x"80",x"31",x"72",x"18",x"10",x"81",x"00",x"00", -- 0x04E8
    x"00",x"00",x"8E",x"84",x"C4",x"BD",x"BA",x"CA", -- 0x04F0
    x"BD",x"BC",x"2F",x"96",x"4F",x"81",x"88",x"25", -- 0x04F8
    x"03",x"7E",x"BB",x"5C",x"BD",x"BC",x"EE",x"96", -- 0x0500
    x"01",x"8B",x"81",x"27",x"F4",x"4A",x"34",x"02", -- 0x0508
    x"8E",x"00",x"40",x"BD",x"B9",x"B9",x"8E",x"84", -- 0x0510
    x"C9",x"BD",x"BE",x"FF",x"0F",x"62",x"35",x"02", -- 0x0518
    x"BD",x"BB",x"48",x"39",x"BD",x"BC",x"6D",x"2B", -- 0x0520
    x"03",x"7E",x"BC",x"EE",x"03",x"54",x"8D",x"F9", -- 0x0528
    x"7E",x"BE",x"E9",x"BD",x"89",x"AE",x"32",x"62", -- 0x0530
    x"86",x"01",x"97",x"D8",x"BD",x"AD",x"01",x"10", -- 0x0538
    x"25",x"29",x"8F",x"BD",x"B7",x"C2",x"1F",x"20", -- 0x0540
    x"83",x"02",x"DE",x"D7",x"D7",x"DC",x"2B",x"BD", -- 0x0548
    x"BD",x"CC",x"BD",x"B9",x"AC",x"8E",x"02",x"DD", -- 0x0550
    x"D6",x"D8",x"26",x"25",x"5F",x"BD",x"86",x"87", -- 0x0558
    x"BD",x"90",x"AA",x"25",x"0B",x"80",x"30",x"34", -- 0x0560
    x"02",x"86",x"0A",x"3D",x"EB",x"E0",x"20",x"ED", -- 0x0568
    x"C0",x"01",x"C9",x"01",x"81",x"41",x"26",x"05", -- 0x0570
    x"BD",x"B9",x"58",x"20",x"BB",x"81",x"4C",x"26", -- 0x0578
    x"0B",x"8D",x"31",x"0F",x"D8",x"BD",x"B9",x"58", -- 0x0580
    x"20",x"C3",x"32",x"62",x"81",x"0D",x"26",x"0D", -- 0x0588
    x"8D",x"22",x"BD",x"B9",x"58",x"8E",x"02",x"DD", -- 0x0590
    x"9F",x"A6",x"7E",x"AC",x"A8",x"81",x"45",x"27", -- 0x0598
    x"F1",x"81",x"51",x"26",x"06",x"BD",x"B9",x"58", -- 0x05A0
    x"7E",x"AC",x"73",x"8D",x"02",x"20",x"AD",x"81", -- 0x05A8
    x"20",x"26",x"10",x"8C",x"C6",x"F9",x"A6",x"84", -- 0x05B0
    x"27",x"08",x"BD",x"A2",x"82",x"30",x"01",x"5A", -- 0x05B8
    x"26",x"F4",x"39",x"81",x"44",x"26",x"48",x"6D", -- 0x05C0
    x"84",x"27",x"F7",x"8D",x"04",x"5A",x"26",x"F7", -- 0x05C8
    x"39",x"0A",x"D7",x"31",x"1F",x"31",x"21",x"A6", -- 0x05D0
    x"21",x"A7",x"A4",x"26",x"F8",x"39",x"81",x"49", -- 0x05D8
    x"27",x"13",x"81",x"58",x"27",x"0D",x"81",x"48", -- 0x05E0
    x"26",x"5C",x"6F",x"84",x"1F",x"10",x"83",x"02", -- 0x05E8
    x"DE",x"D7",x"D7",x"8D",x"BF",x"BD",x"86",x"87", -- 0x05F0
    x"81",x"0D",x"27",x"8E",x"81",x"1B",x"27",x"25", -- 0x05F8
    x"81",x"08",x"26",x"22",x"8C",x"02",x"DD",x"27", -- 0x0600
    x"EC",x"8D",x"45",x"8D",x"C4",x"20",x"E6",x"81", -- 0x0608
    x"43",x"26",x"CB",x"6D",x"84",x"27",x"0E",x"BD", -- 0x0610
    x"86",x"87",x"25",x"02",x"20",x"F5",x"A7",x"80", -- 0x0618
    x"8D",x"37",x"5A",x"26",x"EE",x"39",x"D6",x"D7", -- 0x0620
    x"C1",x"F9",x"26",x"02",x"20",x"C7",x"34",x"10", -- 0x0628
    x"6D",x"80",x"26",x"FC",x"E6",x"82",x"E7",x"01", -- 0x0630
    x"AC",x"E4",x"26",x"F8",x"32",x"62",x"A7",x"80", -- 0x0638
    x"8D",x"17",x"0C",x"D7",x"20",x"AF",x"81",x"08", -- 0x0640
    x"26",x"12",x"8D",x"04",x"5A",x"26",x"FB",x"39", -- 0x0648
    x"8C",x"02",x"DD",x"27",x"D0",x"30",x"1F",x"86", -- 0x0650
    x"08",x"7E",x"A2",x"82",x"81",x"4B",x"27",x"05", -- 0x0658
    x"80",x"53",x"27",x"01",x"39",x"34",x"02",x"8D", -- 0x0660
    x"1E",x"34",x"02",x"A6",x"84",x"27",x"16",x"6D", -- 0x0668
    x"61",x"26",x"06",x"8D",x"E4",x"30",x"01",x"20", -- 0x0670
    x"03",x"BD",x"85",x"D1",x"A6",x"84",x"A1",x"E4", -- 0x0678
    x"26",x"E9",x"5A",x"26",x"E6",x"35",x"A0",x"BD", -- 0x0680
    x"A1",x"71",x"81",x"7F",x"24",x"F9",x"81",x"5F", -- 0x0688
    x"26",x"02",x"86",x"1B",x"81",x"0D",x"27",x"0E", -- 0x0690
    x"81",x"1B",x"27",x"0A",x"81",x"08",x"27",x"06", -- 0x0698
    x"81",x"20",x"25",x"E3",x"1A",x"01",x"39",x"86", -- 0x06A0
    x"4F",x"97",x"AF",x"39",x"96",x"6F",x"34",x"02", -- 0x06A8
    x"BD",x"A5",x"AE",x"BD",x"A4",x"06",x"BD",x"A3", -- 0x06B0
    x"5F",x"D6",x"6C",x"7E",x"A5",x"E4",x"BD",x"B2", -- 0x06B8
    x"6A",x"DC",x"1F",x"34",x"06",x"BD",x"B3",x"57", -- 0x06C0
    x"BD",x"B2",x"67",x"35",x"06",x"1E",x"10",x"9C", -- 0x06C8
    x"1F",x"26",x"51",x"7E",x"B4",x"F4",x"9D",x"9F", -- 0x06D0
    x"BD",x"B2",x"6A",x"BD",x"B3",x"57",x"34",x"10", -- 0x06D8
    x"EC",x"02",x"10",x"93",x"21",x"23",x"04",x"93", -- 0x06E0
    x"27",x"23",x"12",x"E6",x"84",x"BD",x"B5",x"6D", -- 0x06E8
    x"34",x"10",x"AE",x"62",x"BD",x"B6",x"43",x"35", -- 0x06F0
    x"50",x"AF",x"42",x"34",x"40",x"BD",x"B7",x"38", -- 0x06F8
    x"34",x"04",x"5D",x"27",x"1F",x"C6",x"FF",x"81", -- 0x0700
    x"29",x"27",x"03",x"BD",x"B7",x"38",x"34",x"04", -- 0x0708
    x"BD",x"B2",x"67",x"C6",x"B3",x"BD",x"B2",x"6F", -- 0x0710
    x"8D",x"2E",x"1F",x"13",x"AE",x"62",x"A6",x"84", -- 0x0718
    x"A0",x"61",x"24",x"03",x"7E",x"B4",x"4A",x"4C", -- 0x0720
    x"A1",x"E4",x"24",x"02",x"A7",x"E4",x"A6",x"61", -- 0x0728
    x"1E",x"89",x"AE",x"02",x"5A",x"3A",x"4D",x"27", -- 0x0730
    x"0D",x"A1",x"E4",x"23",x"02",x"A6",x"E4",x"1F", -- 0x0738
    x"89",x"1E",x"31",x"BD",x"A5",x"9A",x"35",x"96", -- 0x0740
    x"BD",x"B1",x"56",x"7E",x"B6",x"54",x"BD",x"B2", -- 0x0748
    x"6A",x"BD",x"B7",x"0B",x"34",x"04",x"BD",x"B2", -- 0x0750
    x"6D",x"BD",x"B1",x"56",x"BD",x"B2",x"67",x"96", -- 0x0758
    x"06",x"26",x"05",x"BD",x"B7",x"0E",x"20",x"03", -- 0x0760
    x"BD",x"B6",x"A4",x"34",x"04",x"E6",x"61",x"BD", -- 0x0768
    x"B5",x"0F",x"35",x"06",x"27",x"05",x"A7",x"80", -- 0x0770
    x"5A",x"26",x"FB",x"7E",x"B6",x"9B",x"BD",x"B2", -- 0x0778
    x"6A",x"BD",x"B1",x"56",x"C6",x"01",x"34",x"04", -- 0x0780
    x"96",x"06",x"26",x"10",x"BD",x"B7",x"0E",x"E7", -- 0x0788
    x"E4",x"27",x"91",x"BD",x"B2",x"6D",x"BD",x"B1", -- 0x0790
    x"56",x"BD",x"B1",x"46",x"9E",x"52",x"34",x"10", -- 0x0798
    x"BD",x"B2",x"6D",x"BD",x"87",x"48",x"34",x"14", -- 0x07A0
    x"BD",x"B2",x"67",x"AE",x"63",x"BD",x"B6",x"59", -- 0x07A8
    x"34",x"04",x"E1",x"66",x"25",x"23",x"A6",x"61", -- 0x07B0
    x"27",x"1C",x"E6",x"66",x"5A",x"3A",x"31",x"84", -- 0x07B8
    x"EE",x"62",x"E6",x"61",x"A6",x"E4",x"A0",x"66", -- 0x07C0
    x"4C",x"A1",x"61",x"25",x"0C",x"A6",x"80",x"A1", -- 0x07C8
    x"C0",x"26",x"0C",x"5A",x"26",x"F7",x"E6",x"66", -- 0x07D0
    x"21",x"5F",x"32",x"67",x"7E",x"B4",x"F3",x"6C", -- 0x07D8
    x"66",x"30",x"21",x"20",x"D9",x"81",x"26",x"26", -- 0x07E0
    x"5C",x"32",x"62",x"0F",x"52",x"0F",x"53",x"8E", -- 0x07E8
    x"00",x"52",x"9D",x"9F",x"81",x"4F",x"27",x"12", -- 0x07F0
    x"81",x"48",x"27",x"23",x"9D",x"A5",x"20",x"0C", -- 0x07F8
    x"81",x"38",x"10",x"22",x"2A",x"71",x"C6",x"03", -- 0x0800
    x"8D",x"2A",x"9D",x"9F",x"25",x"F2",x"0F",x"50", -- 0x0808
    x"0F",x"51",x"0F",x"06",x"0F",x"63",x"0F",x"54", -- 0x0810
    x"C6",x"A0",x"D7",x"4F",x"7E",x"BA",x"1C",x"9D", -- 0x0818
    x"9F",x"25",x"0B",x"BD",x"B3",x"A2",x"25",x"E6", -- 0x0820
    x"81",x"47",x"24",x"E2",x"80",x"07",x"C6",x"04", -- 0x0828
    x"8D",x"02",x"20",x"EB",x"68",x"01",x"69",x"84", -- 0x0830
    x"10",x"25",x"32",x"56",x"5A",x"26",x"F5",x"80", -- 0x0838
    x"30",x"AB",x"01",x"A7",x"01",x"39",x"35",x"40", -- 0x0840
    x"0F",x"06",x"9E",x"A6",x"9D",x"9F",x"81",x"26", -- 0x0848
    x"27",x"99",x"81",x"CC",x"27",x"5E",x"81",x"FF", -- 0x0850
    x"26",x"08",x"9D",x"9F",x"81",x"83",x"10",x"27", -- 0x0858
    x"00",x"CA",x"9F",x"A6",x"6E",x"C4",x"9E",x"68", -- 0x0860
    x"30",x"01",x"26",x"D9",x"C6",x"16",x"7E",x"AC", -- 0x0868
    x"46",x"AE",x"9F",x"00",x"A6",x"8C",x"FF",x"83", -- 0x0870
    x"10",x"27",x"00",x"93",x"8D",x"23",x"8D",x"E6", -- 0x0878
    x"BD",x"B2",x"6A",x"C6",x"80",x"D7",x"08",x"BD", -- 0x0880
    x"B3",x"57",x"8D",x"25",x"BD",x"B2",x"67",x"C6", -- 0x0888
    x"B3",x"BD",x"B2",x"6F",x"9E",x"4B",x"DC",x"A6", -- 0x0890
    x"ED",x"84",x"DC",x"39",x"ED",x"02",x"7E",x"AE", -- 0x0898
    x"E0",x"C6",x"CC",x"BD",x"B2",x"6F",x"C6",x"80", -- 0x08A0
    x"D7",x"08",x"8A",x"80",x"BD",x"B3",x"5C",x"9F", -- 0x08A8
    x"4B",x"7E",x"B1",x"43",x"8D",x"EB",x"34",x"10", -- 0x08B0
    x"BD",x"B2",x"62",x"8D",x"F4",x"35",x"40",x"C6", -- 0x08B8
    x"32",x"AE",x"42",x"27",x"A9",x"10",x"9E",x"A6", -- 0x08C0
    x"EE",x"C4",x"DF",x"A6",x"A6",x"04",x"34",x"02", -- 0x08C8
    x"EC",x"84",x"EE",x"02",x"34",x"76",x"BD",x"BC", -- 0x08D0
    x"35",x"BD",x"B1",x"41",x"35",x"76",x"ED",x"84", -- 0x08D8
    x"EF",x"02",x"35",x"02",x"A7",x"04",x"9D",x"A5", -- 0x08E0
    x"10",x"26",x"29",x"8B",x"10",x"9F",x"A6",x"39", -- 0x08E8
    x"C1",x"32",x"25",x"FB",x"BD",x"A7",x"E9",x"BD", -- 0x08F0
    x"A9",x"74",x"BD",x"AD",x"33",x"0F",x"6F",x"BD", -- 0x08F8
    x"B9",x"5C",x"BD",x"B9",x"AF",x"8E",x"88",x"D9", -- 0x0900
    x"7E",x"AC",x"60",x"55",x"46",x"4E",x"45",x"9D", -- 0x0908
    x"9F",x"8D",x"09",x"34",x"10",x"8D",x"2D",x"35", -- 0x0910
    x"40",x"AF",x"C4",x"39",x"5F",x"9D",x"9F",x"24", -- 0x0918
    x"06",x"80",x"30",x"1F",x"89",x"9D",x"9F",x"9E", -- 0x0920
    x"B0",x"58",x"3A",x"39",x"8D",x"EE",x"AE",x"84", -- 0x0928
    x"34",x"10",x"BD",x"B2",x"62",x"8E",x"00",x"4F", -- 0x0930
    x"96",x"06",x"27",x"07",x"BD",x"B6",x"57",x"9E", -- 0x0938
    x"52",x"96",x"06",x"39",x"C6",x"B3",x"BD",x"B2", -- 0x0940
    x"6F",x"7E",x"B7",x"3D",x"B6",x"FF",x"03",x"2B", -- 0x0948
    x"01",x"3B",x"B6",x"FF",x"02",x"BE",x"01",x"12", -- 0x0950
    x"30",x"01",x"BF",x"01",x"12",x"7E",x"9C",x"3E", -- 0x0958
    x"9D",x"9F",x"8D",x"E0",x"BF",x"01",x"12",x"39", -- 0x0960
    x"BE",x"01",x"12",x"9F",x"52",x"7E",x"88",x"0E", -- 0x0968
    x"10",x"27",x"2A",x"D6",x"BD",x"AF",x"67",x"BD", -- 0x0970
    x"AD",x"01",x"9F",x"D3",x"9D",x"A5",x"27",x"10", -- 0x0978
    x"81",x"AC",x"26",x"3B",x"9D",x"9F",x"27",x"04", -- 0x0980
    x"8D",x"24",x"20",x"04",x"86",x"FF",x"97",x"2B", -- 0x0988
    x"DE",x"D3",x"8C",x"EE",x"C4",x"EC",x"C4",x"27", -- 0x0990
    x"06",x"EC",x"42",x"93",x"2B",x"23",x"F4",x"9E", -- 0x0998
    x"D3",x"8D",x"15",x"BD",x"AD",x"21",x"9E",x"D3", -- 0x09A0
    x"BD",x"AC",x"F1",x"7E",x"AC",x"73",x"BD",x"AF", -- 0x09A8
    x"67",x"7E",x"A5",x"C7",x"A6",x"C0",x"A7",x"80", -- 0x09B0
    x"11",x"93",x"1B",x"26",x"F7",x"9F",x"1B",x"39", -- 0x09B8
    x"BD",x"88",x"66",x"9D",x"9F",x"81",x"23",x"26", -- 0x09C0
    x"09",x"BD",x"A5",x"A5",x"BD",x"A3",x"ED",x"BD", -- 0x09C8
    x"B2",x"6D",x"81",x"22",x"26",x"0B",x"BD",x"B2", -- 0x09D0
    x"44",x"C6",x"3B",x"BD",x"B2",x"6F",x"BD",x"B9", -- 0x09D8
    x"9F",x"32",x"7E",x"BD",x"B0",x"35",x"32",x"62", -- 0x09E0
    x"0F",x"6F",x"BD",x"B3",x"57",x"9F",x"3B",x"BD", -- 0x09E8
    x"B1",x"46",x"8E",x"02",x"DC",x"4F",x"BD",x"B5", -- 0x09F0
    x"1A",x"7E",x"AF",x"A4",x"BD",x"AF",x"67",x"9E", -- 0x09F8
    x"2B",x"39",x"9E",x"D1",x"9F",x"2B",x"7E",x"AD", -- 0x0A00
    x"01",x"BD",x"AD",x"26",x"CC",x"00",x"0A",x"DD", -- 0x0A08
    x"D5",x"DD",x"CF",x"5F",x"DD",x"D1",x"9D",x"A5", -- 0x0A10
    x"24",x"06",x"8D",x"E0",x"9F",x"D5",x"9D",x"A5", -- 0x0A18
    x"27",x"1B",x"BD",x"B2",x"6D",x"24",x"06",x"8D", -- 0x0A20
    x"D3",x"9F",x"D1",x"9D",x"A5",x"27",x"0E",x"BD", -- 0x0A28
    x"B2",x"6D",x"24",x"06",x"8D",x"C6",x"9F",x"CF", -- 0x0A30
    x"27",x"49",x"BD",x"A5",x"C7",x"8D",x"C3",x"9F", -- 0x0A38
    x"D3",x"9E",x"D5",x"8D",x"BF",x"9C",x"D3",x"25", -- 0x0A40
    x"3A",x"8D",x"1C",x"BD",x"8A",x"DD",x"BD",x"AC", -- 0x0A48
    x"EF",x"8D",x"AF",x"9F",x"D3",x"8D",x"3A",x"8D", -- 0x0A50
    x"0F",x"8D",x"36",x"BD",x"8B",x"7B",x"BD",x"AD", -- 0x0A58
    x"26",x"BD",x"AC",x"EF",x"7E",x"AC",x"73",x"86", -- 0x0A60
    x"4F",x"97",x"D8",x"9E",x"D3",x"DC",x"D5",x"8D", -- 0x0A68
    x"15",x"0D",x"D8",x"26",x"02",x"ED",x"02",x"AE", -- 0x0A70
    x"84",x"8D",x"0B",x"D3",x"CF",x"25",x"04",x"81", -- 0x0A78
    x"FA",x"25",x"EE",x"7E",x"B4",x"4A",x"34",x"06", -- 0x0A80
    x"EC",x"84",x"35",x"06",x"26",x"02",x"32",x"62", -- 0x0A88
    x"39",x"9E",x"19",x"30",x"1F",x"30",x"01",x"8D", -- 0x0A90
    x"ED",x"30",x"03",x"30",x"01",x"A6",x"84",x"27", -- 0x0A98
    x"F4",x"9F",x"0F",x"4A",x"27",x"0C",x"4A",x"27", -- 0x0AA0
    x"2A",x"4A",x"26",x"EF",x"86",x"03",x"A7",x"80", -- 0x0AA8
    x"20",x"E7",x"EC",x"01",x"6A",x"02",x"27",x"01", -- 0x0AB0
    x"4F",x"E6",x"03",x"6A",x"04",x"27",x"01",x"5F", -- 0x0AB8
    x"ED",x"01",x"DD",x"2B",x"BD",x"AD",x"01",x"9E", -- 0x0AC0
    x"0F",x"25",x"E1",x"DC",x"47",x"6C",x"80",x"ED", -- 0x0AC8
    x"84",x"20",x"C6",x"6F",x"84",x"AE",x"01",x"AE", -- 0x0AD0
    x"02",x"9F",x"47",x"20",x"EA",x"9E",x"19",x"20", -- 0x0AD8
    x"04",x"9E",x"A6",x"30",x"01",x"8D",x"9F",x"30", -- 0x0AE0
    x"02",x"30",x"01",x"9F",x"A6",x"9D",x"9F",x"4D", -- 0x0AE8
    x"27",x"EF",x"2A",x"F9",x"9E",x"A6",x"81",x"FF", -- 0x0AF0
    x"27",x"EF",x"BD",x"01",x"A0",x"81",x"A7",x"27", -- 0x0AF8
    x"12",x"81",x"84",x"27",x"0E",x"81",x"81",x"26", -- 0x0B00
    x"E4",x"9D",x"9F",x"81",x"A5",x"27",x"04",x"81", -- 0x0B08
    x"A6",x"26",x"D8",x"9D",x"9F",x"25",x"04",x"9D", -- 0x0B10
    x"A5",x"20",x"D4",x"9E",x"A6",x"34",x"10",x"BD", -- 0x0B18
    x"AF",x"67",x"9E",x"A6",x"A6",x"82",x"BD",x"90", -- 0x0B20
    x"AA",x"25",x"F9",x"30",x"01",x"1F",x"10",x"E0", -- 0x0B28
    x"61",x"C0",x"05",x"27",x"20",x"25",x"0A",x"33", -- 0x0B30
    x"84",x"50",x"30",x"85",x"BD",x"89",x"B8",x"20", -- 0x0B38
    x"14",x"9F",x"47",x"9E",x"1B",x"9F",x"43",x"50", -- 0x0B40
    x"30",x"85",x"9F",x"41",x"9F",x"1B",x"BD",x"AC", -- 0x0B48
    x"1E",x"9E",x"45",x"9F",x"A6",x"35",x"10",x"86", -- 0x0B50
    x"01",x"A7",x"84",x"A7",x"02",x"A7",x"04",x"D6", -- 0x0B58
    x"2B",x"26",x"04",x"C6",x"01",x"6C",x"02",x"E7", -- 0x0B60
    x"01",x"D6",x"2C",x"26",x"04",x"C6",x"01",x"6C", -- 0x0B68
    x"04",x"E7",x"03",x"9D",x"A5",x"81",x"2C",x"27", -- 0x0B70
    x"9A",x"20",x"9C",x"9E",x"19",x"30",x"1F",x"30", -- 0x0B78
    x"01",x"EC",x"02",x"DD",x"68",x"BD",x"8A",x"86", -- 0x0B80
    x"30",x"03",x"30",x"01",x"A6",x"84",x"27",x"EF", -- 0x0B88
    x"4A",x"27",x"1B",x"80",x"02",x"26",x"F3",x"34", -- 0x0B90
    x"10",x"8E",x"8B",x"D8",x"BD",x"B9",x"9C",x"AE", -- 0x0B98
    x"E4",x"EC",x"01",x"BD",x"BD",x"CC",x"BD",x"BD", -- 0x0BA0
    x"C5",x"BD",x"B9",x"58",x"35",x"10",x"34",x"10", -- 0x0BA8
    x"EC",x"01",x"DD",x"52",x"BD",x"88",x"0E",x"BD", -- 0x0BB0
    x"BD",x"D9",x"35",x"40",x"C6",x"05",x"30",x"01", -- 0x0BB8
    x"A6",x"84",x"27",x"05",x"5A",x"A7",x"C0",x"20", -- 0x0BC0
    x"F5",x"30",x"C4",x"5D",x"27",x"BE",x"31",x"C4", -- 0x0BC8
    x"33",x"C5",x"BD",x"89",x"B8",x"30",x"A4",x"20", -- 0x0BD0
    x"B3",x"55",x"4C",x"20",x"00",x"BD",x"B7",x"40", -- 0x0BD8
    x"8E",x"03",x"D9",x"C6",x"04",x"34",x"04",x"5F", -- 0x0BE0
    x"86",x"04",x"08",x"53",x"09",x"52",x"59",x"4A", -- 0x0BE8
    x"26",x"F8",x"5D",x"26",x"0A",x"A6",x"E4",x"4A", -- 0x0BF0
    x"27",x"05",x"8C",x"03",x"D9",x"27",x"0C",x"CB", -- 0x0BF8
    x"30",x"C1",x"39",x"23",x"02",x"CB",x"07",x"E7", -- 0x0C00
    x"80",x"6F",x"84",x"35",x"04",x"5A",x"26",x"D5", -- 0x0C08
    x"32",x"62",x"8E",x"03",x"D8",x"7E",x"B5",x"18", -- 0x0C10
    x"BD",x"A4",x"29",x"1A",x"50",x"86",x"0A",x"B7", -- 0x0C18
    x"FF",x"90",x"7F",x"FF",x"DE",x"7E",x"C0",x"00", -- 0x0C20
    x"7F",x"FE",x"ED",x"7F",x"FF",x"23",x"86",x"CC", -- 0x0C28
    x"B7",x"FF",x"90",x"7F",x"FF",x"DE",x"39",x"34", -- 0x0C30
    x"16",x"9E",x"88",x"D6",x"E7",x"10",x"26",x"6B", -- 0x0C38
    x"6D",x"E6",x"61",x"7E",x"A3",x"0E",x"34",x"01", -- 0x0C40
    x"0D",x"E7",x"27",x"03",x"7E",x"F6",x"AD",x"35", -- 0x0C48
    x"01",x"7E",x"A9",x"13",x"12",x"C7",x"5D",x"27", -- 0x0C50
    x"06",x"BD",x"AD",x"19",x"7E",x"AC",x"7C",x"7E", -- 0x0C58
    x"A6",x"16",x"9D",x"9F",x"81",x"4D",x"10",x"26", -- 0x0C60
    x"18",x"2E",x"0F",x"78",x"9D",x"9F",x"BD",x"A5", -- 0x0C68
    x"78",x"BD",x"A6",x"48",x"7D",x"01",x"E4",x"10", -- 0x0C70
    x"27",x"18",x"8A",x"FE",x"01",x"E2",x"0A",x"6F", -- 0x0C78
    x"BD",x"A6",x"35",x"1F",x"30",x"83",x"02",x"00", -- 0x0C80
    x"26",x"D5",x"9E",x"8A",x"9D",x"A5",x"27",x"06", -- 0x0C88
    x"BD",x"B2",x"6D",x"BD",x"B7",x"3D",x"9F",x"D3", -- 0x0C90
    x"BD",x"A5",x"C7",x"8D",x"29",x"34",x"02",x"8D", -- 0x0C98
    x"1E",x"1F",x"02",x"8D",x"1A",x"D3",x"D3",x"DD", -- 0x0CA0
    x"9D",x"1F",x"01",x"A6",x"E0",x"10",x"26",x"17", -- 0x0CA8
    x"7C",x"8D",x"13",x"A7",x"84",x"A1",x"80",x"26", -- 0x0CB0
    x"14",x"31",x"3F",x"26",x"F4",x"20",x"DC",x"8D", -- 0x0CB8
    x"00",x"8D",x"03",x"1E",x"89",x"39",x"BD",x"A1", -- 0x0CC0
    x"76",x"0D",x"70",x"27",x"F8",x"7E",x"A6",x"19", -- 0x0CC8
    x"8D",x"42",x"34",x"06",x"4C",x"27",x"06",x"DE", -- 0x0CD0
    x"8A",x"8D",x"09",x"35",x"86",x"C6",x"34",x"7E", -- 0x0CD8
    x"AC",x"46",x"DE",x"7E",x"30",x"41",x"9F",x"7E", -- 0x0CE0
    x"8E",x"01",x"DA",x"BD",x"8D",x"7C",x"7E",x"A6", -- 0x0CE8
    x"44",x"96",x"6F",x"81",x"FD",x"26",x"0A",x"32", -- 0x0CF0
    x"62",x"0F",x"70",x"0D",x"79",x"26",x"03",x"03", -- 0x0CF8
    x"70",x"39",x"34",x"74",x"9E",x"7A",x"A6",x"80", -- 0x0D00
    x"34",x"02",x"9F",x"7A",x"0A",x"79",x"26",x"02", -- 0x0D08
    x"8D",x"D0",x"35",x"F6",x"4F",x"34",x"16",x"31", -- 0x0D10
    x"E4",x"20",x"02",x"8D",x"2B",x"86",x"8A",x"8D", -- 0x0D18
    x"37",x"26",x"F8",x"8E",x"01",x"D2",x"A6",x"80", -- 0x0D20
    x"BD",x"8E",x"04",x"8C",x"01",x"DA",x"26",x"F6", -- 0x0D28
    x"8D",x"30",x"26",x"E7",x"8D",x"3C",x"26",x"E3", -- 0x0D30
    x"A7",x"22",x"8D",x"36",x"26",x"DD",x"A7",x"23", -- 0x0D38
    x"8D",x"29",x"26",x"D7",x"32",x"62",x"35",x"86", -- 0x0D40
    x"6C",x"A4",x"A6",x"A4",x"81",x"05",x"25",x"1A", -- 0x0D48
    x"86",x"BC",x"BD",x"8E",x"0C",x"7E",x"A6",x"19", -- 0x0D50
    x"34",x"02",x"8D",x"5C",x"26",x"02",x"A1",x"E4", -- 0x0D58
    x"35",x"82",x"A6",x"21",x"8D",x"52",x"26",x"02", -- 0x0D60
    x"81",x"C8",x"39",x"8D",x"05",x"26",x"FB",x"A6", -- 0x0D68
    x"21",x"39",x"8D",x"48",x"34",x"03",x"A8",x"21", -- 0x0D70
    x"A7",x"21",x"35",x"83",x"4F",x"34",x"76",x"68", -- 0x0D78
    x"67",x"69",x"66",x"64",x"67",x"31",x"E4",x"20", -- 0x0D80
    x"02",x"8D",x"BD",x"86",x"97",x"8D",x"C9",x"26", -- 0x0D88
    x"F8",x"A6",x"26",x"8D",x"6F",x"A6",x"27",x"8D", -- 0x0D90
    x"6B",x"8D",x"C7",x"26",x"EC",x"8D",x"D3",x"26", -- 0x0D98
    x"E8",x"A7",x"24",x"AE",x"22",x"C6",x"80",x"8D", -- 0x0DA0
    x"C9",x"26",x"DE",x"A7",x"80",x"5A",x"26",x"F7", -- 0x0DA8
    x"8D",x"B9",x"26",x"D5",x"32",x"64",x"35",x"96", -- 0x0DB0
    x"6F",x"21",x"8D",x"50",x"4F",x"34",x"15",x"1A", -- 0x0DB8
    x"50",x"96",x"E7",x"9E",x"8A",x"8D",x"1F",x"24", -- 0x0DC0
    x"FC",x"8D",x"1B",x"25",x"FC",x"8D",x"2A",x"C6", -- 0x0DC8
    x"01",x"34",x"04",x"4F",x"8D",x"21",x"F6",x"FF", -- 0x0DD0
    x"22",x"56",x"24",x"02",x"AA",x"E4",x"68",x"E4", -- 0x0DD8
    x"24",x"F2",x"32",x"61",x"35",x"95",x"F6",x"FF", -- 0x0DE0
    x"22",x"56",x"30",x"01",x"26",x"08",x"4A",x"26", -- 0x0DE8
    x"05",x"32",x"62",x"35",x"15",x"4C",x"39",x"8D", -- 0x0DF0
    x"00",x"34",x"02",x"96",x"E6",x"21",x"FE",x"4A", -- 0x0DF8
    x"26",x"FB",x"35",x"82",x"34",x"02",x"A8",x"21", -- 0x0E00
    x"A7",x"21",x"35",x"02",x"34",x"07",x"1A",x"50", -- 0x0E08
    x"8D",x"E5",x"8D",x"E3",x"7F",x"FF",x"20",x"8D", -- 0x0E10
    x"DE",x"C6",x"01",x"34",x"04",x"A6",x"62",x"A4", -- 0x0E18
    x"E4",x"27",x"02",x"86",x"02",x"B7",x"FF",x"20", -- 0x0E20
    x"8D",x"CD",x"68",x"E4",x"24",x"EF",x"86",x"02", -- 0x0E28
    x"B7",x"FF",x"20",x"32",x"61",x"35",x"87",x"86", -- 0x0E30
    x"01",x"97",x"D9",x"5A",x"BD",x"8F",x"D8",x"9D", -- 0x0E38
    x"A5",x"10",x"27",x"00",x"93",x"D7",x"D3",x"BD", -- 0x0E40
    x"B1",x"56",x"BD",x"B1",x"46",x"9E",x"52",x"9F", -- 0x0E48
    x"4D",x"D6",x"D9",x"BD",x"B6",x"AD",x"BD",x"B9", -- 0x0E50
    x"9F",x"9E",x"52",x"D6",x"D9",x"E0",x"84",x"5A", -- 0x0E58
    x"10",x"2B",x"01",x"4F",x"BD",x"B9",x"AC",x"20", -- 0x0E60
    x"F6",x"D7",x"D3",x"9F",x"0F",x"86",x"02",x"97", -- 0x0E68
    x"D9",x"A6",x"84",x"81",x"25",x"27",x"C4",x"81", -- 0x0E70
    x"20",x"26",x"07",x"0C",x"D9",x"30",x"01",x"5A", -- 0x0E78
    x"26",x"EF",x"9E",x"0F",x"D6",x"D3",x"86",x"25", -- 0x0E80
    x"BD",x"8F",x"D8",x"BD",x"A2",x"82",x"20",x"29", -- 0x0E88
    x"81",x"CD",x"27",x"01",x"39",x"32",x"62",x"BD", -- 0x0E90
    x"B1",x"58",x"BD",x"B1",x"46",x"C6",x"3B",x"BD", -- 0x0E98
    x"B2",x"6F",x"9E",x"52",x"9F",x"D5",x"20",x"06", -- 0x0EA0
    x"96",x"D7",x"27",x"08",x"9E",x"D5",x"0F",x"D7", -- 0x0EA8
    x"E6",x"84",x"26",x"03",x"7E",x"B4",x"4A",x"AE", -- 0x0EB0
    x"02",x"0F",x"DA",x"0F",x"D9",x"A6",x"80",x"81", -- 0x0EB8
    x"21",x"10",x"27",x"FF",x"72",x"81",x"23",x"27", -- 0x0EC0
    x"5B",x"5A",x"26",x"16",x"BD",x"8F",x"D8",x"BD", -- 0x0EC8
    x"A2",x"82",x"9D",x"A5",x"26",x"D2",x"96",x"D7", -- 0x0ED0
    x"26",x"03",x"BD",x"B9",x"58",x"9E",x"D5",x"7E", -- 0x0ED8
    x"B6",x"59",x"81",x"2B",x"26",x"09",x"BD",x"8F", -- 0x0EE0
    x"D8",x"86",x"08",x"97",x"DA",x"20",x"CC",x"81", -- 0x0EE8
    x"2E",x"27",x"4E",x"81",x"25",x"10",x"27",x"FF", -- 0x0EF0
    x"70",x"A1",x"84",x"26",x"8B",x"81",x"24",x"27", -- 0x0EF8
    x"19",x"81",x"2A",x"26",x"F6",x"96",x"DA",x"8A", -- 0x0F00
    x"20",x"97",x"DA",x"C1",x"02",x"25",x"11",x"A6", -- 0x0F08
    x"01",x"81",x"24",x"26",x"0B",x"5A",x"30",x"01", -- 0x0F10
    x"0C",x"D9",x"96",x"DA",x"8A",x"10",x"97",x"DA", -- 0x0F18
    x"30",x"01",x"0C",x"D9",x"0F",x"D8",x"0C",x"D9", -- 0x0F20
    x"5A",x"27",x"49",x"A6",x"80",x"81",x"2E",x"27", -- 0x0F28
    x"1E",x"81",x"23",x"27",x"F1",x"81",x"2C",x"26", -- 0x0F30
    x"21",x"96",x"DA",x"8A",x"40",x"97",x"DA",x"20", -- 0x0F38
    x"E5",x"A6",x"84",x"81",x"23",x"10",x"26",x"FF", -- 0x0F40
    x"3F",x"86",x"01",x"97",x"D8",x"30",x"01",x"0C", -- 0x0F48
    x"D8",x"5A",x"27",x"20",x"A6",x"80",x"81",x"23", -- 0x0F50
    x"27",x"F5",x"81",x"5E",x"26",x"16",x"A1",x"84", -- 0x0F58
    x"26",x"12",x"A1",x"01",x"26",x"0E",x"A1",x"02", -- 0x0F60
    x"26",x"0A",x"C1",x"04",x"25",x"06",x"C0",x"04", -- 0x0F68
    x"30",x"04",x"0C",x"DA",x"30",x"1F",x"0C",x"D9", -- 0x0F70
    x"96",x"DA",x"85",x"08",x"26",x"18",x"0A",x"D9", -- 0x0F78
    x"5D",x"27",x"13",x"A6",x"84",x"80",x"2D",x"27", -- 0x0F80
    x"06",x"81",x"FE",x"26",x"09",x"86",x"08",x"8A", -- 0x0F88
    x"04",x"9A",x"DA",x"97",x"DA",x"5A",x"9D",x"A5", -- 0x0F90
    x"10",x"27",x"FF",x"3C",x"D7",x"D3",x"BD",x"B1", -- 0x0F98
    x"41",x"96",x"D9",x"9B",x"D8",x"81",x"11",x"10", -- 0x0FA0
    x"22",x"24",x"9F",x"BD",x"8F",x"E5",x"30",x"1F", -- 0x0FA8
    x"BD",x"B9",x"9C",x"0F",x"D7",x"9D",x"A5",x"27", -- 0x0FB0
    x"0D",x"97",x"D7",x"81",x"3B",x"27",x"05",x"BD", -- 0x0FB8
    x"B2",x"6D",x"20",x"02",x"9D",x"9F",x"9E",x"D5", -- 0x0FC0
    x"E6",x"84",x"D0",x"D3",x"AE",x"02",x"3A",x"D6", -- 0x0FC8
    x"D3",x"10",x"26",x"FE",x"E4",x"7E",x"8E",x"D2", -- 0x0FD0
    x"34",x"02",x"86",x"2B",x"0D",x"DA",x"27",x"03", -- 0x0FD8
    x"BD",x"A2",x"82",x"35",x"82",x"CE",x"03",x"DB", -- 0x0FE0
    x"C6",x"20",x"96",x"DA",x"85",x"08",x"27",x"02", -- 0x0FE8
    x"C6",x"2B",x"0D",x"54",x"2A",x"04",x"0F",x"54", -- 0x0FF0
    x"C6",x"2D",x"E7",x"C0",x"C6",x"30",x"E7",x"C0", -- 0x0FF8
    x"84",x"01",x"10",x"26",x"01",x"07",x"8E",x"BD", -- 0x1000
    x"C0",x"BD",x"BC",x"A0",x"2B",x"15",x"BD",x"BD", -- 0x1008
    x"D9",x"A6",x"80",x"26",x"FC",x"A6",x"82",x"A7", -- 0x1010
    x"01",x"8C",x"03",x"DA",x"26",x"F7",x"86",x"25", -- 0x1018
    x"A7",x"84",x"39",x"96",x"4F",x"97",x"47",x"27", -- 0x1020
    x"03",x"BD",x"91",x"CD",x"96",x"47",x"10",x"2B", -- 0x1028
    x"00",x"81",x"40",x"9B",x"D9",x"80",x"09",x"BD", -- 0x1030
    x"90",x"EA",x"BD",x"92",x"63",x"BD",x"92",x"02", -- 0x1038
    x"96",x"47",x"BD",x"92",x"81",x"96",x"47",x"BD", -- 0x1040
    x"92",x"49",x"96",x"D8",x"26",x"02",x"33",x"5F", -- 0x1048
    x"4A",x"BD",x"90",x"EA",x"BD",x"91",x"85",x"4D", -- 0x1050
    x"27",x"06",x"C1",x"2A",x"27",x"02",x"E7",x"C0", -- 0x1058
    x"6F",x"C4",x"8E",x"03",x"DA",x"30",x"01",x"9F", -- 0x1060
    x"0F",x"96",x"3A",x"90",x"10",x"90",x"D9",x"27", -- 0x1068
    x"38",x"A6",x"84",x"81",x"20",x"27",x"EE",x"81", -- 0x1070
    x"2A",x"27",x"EA",x"4F",x"34",x"02",x"A6",x"80", -- 0x1078
    x"81",x"2D",x"27",x"F8",x"81",x"2B",x"27",x"F4", -- 0x1080
    x"81",x"24",x"27",x"F0",x"81",x"30",x"26",x"0E", -- 0x1088
    x"A6",x"01",x"8D",x"16",x"25",x"08",x"35",x"02", -- 0x1090
    x"A7",x"82",x"26",x"FA",x"20",x"C7",x"35",x"02", -- 0x1098
    x"4D",x"26",x"FB",x"9E",x"0F",x"86",x"25",x"A7", -- 0x10A0
    x"82",x"39",x"81",x"30",x"25",x"04",x"80",x"3A", -- 0x10A8
    x"80",x"C6",x"39",x"96",x"D8",x"27",x"01",x"4A", -- 0x10B0
    x"9B",x"47",x"2B",x"01",x"4F",x"34",x"02",x"2A", -- 0x10B8
    x"0A",x"34",x"02",x"BD",x"BB",x"82",x"35",x"02", -- 0x10C0
    x"4C",x"20",x"F4",x"96",x"47",x"A0",x"E0",x"97", -- 0x10C8
    x"47",x"8B",x"09",x"2B",x"19",x"96",x"D9",x"80", -- 0x10D0
    x"09",x"90",x"47",x"8D",x"0D",x"BD",x"92",x"63", -- 0x10D8
    x"20",x"1D",x"34",x"02",x"86",x"30",x"A7",x"C0", -- 0x10E0
    x"35",x"02",x"4A",x"2A",x"F5",x"39",x"96",x"D9", -- 0x10E8
    x"8D",x"F8",x"BD",x"92",x"4D",x"86",x"F7",x"90", -- 0x10F0
    x"47",x"8D",x"EF",x"0F",x"45",x"0F",x"D7",x"BD", -- 0x10F8
    x"92",x"02",x"96",x"D8",x"26",x"02",x"DE",x"39", -- 0x1100
    x"9B",x"47",x"16",x"FF",x"43",x"96",x"4F",x"34", -- 0x1108
    x"02",x"27",x"03",x"BD",x"91",x"CD",x"96",x"D8", -- 0x1110
    x"27",x"01",x"4A",x"9B",x"D9",x"7F",x"03",x"DA", -- 0x1118
    x"D6",x"DA",x"C4",x"04",x"26",x"03",x"73",x"03", -- 0x1120
    x"DA",x"BB",x"03",x"DA",x"80",x"09",x"34",x"02", -- 0x1128
    x"2A",x"0A",x"34",x"02",x"BD",x"BB",x"82",x"35", -- 0x1130
    x"02",x"4C",x"20",x"F4",x"A6",x"E4",x"2B",x"01", -- 0x1138
    x"4F",x"40",x"9B",x"D9",x"4C",x"BB",x"03",x"DA", -- 0x1140
    x"97",x"45",x"0F",x"D7",x"BD",x"92",x"02",x"35", -- 0x1148
    x"02",x"BD",x"92",x"81",x"96",x"D8",x"26",x"02", -- 0x1150
    x"33",x"5F",x"E6",x"E0",x"27",x"09",x"D6",x"47", -- 0x1158
    x"CB",x"09",x"D0",x"D9",x"F0",x"03",x"DA",x"86", -- 0x1160
    x"2B",x"5D",x"2A",x"03",x"86",x"2D",x"50",x"A7", -- 0x1168
    x"41",x"86",x"45",x"A7",x"C1",x"86",x"2F",x"4C", -- 0x1170
    x"C0",x"0A",x"24",x"FB",x"CB",x"3A",x"ED",x"C1", -- 0x1178
    x"6F",x"C4",x"7E",x"90",x"54",x"8E",x"03",x"DB", -- 0x1180
    x"E6",x"84",x"34",x"04",x"86",x"20",x"D6",x"DA", -- 0x1188
    x"C5",x"20",x"35",x"04",x"27",x"08",x"86",x"2A", -- 0x1190
    x"C1",x"20",x"26",x"02",x"1F",x"89",x"34",x"04", -- 0x1198
    x"A7",x"80",x"E6",x"84",x"27",x"10",x"C1",x"45", -- 0x11A0
    x"27",x"0C",x"C1",x"30",x"27",x"F2",x"C1",x"2C", -- 0x11A8
    x"27",x"EE",x"C1",x"2E",x"26",x"04",x"86",x"30", -- 0x11B0
    x"A7",x"82",x"96",x"DA",x"85",x"10",x"27",x"04", -- 0x11B8
    x"C6",x"24",x"E7",x"82",x"84",x"04",x"35",x"04", -- 0x11C0
    x"26",x"02",x"E7",x"82",x"39",x"34",x"40",x"4F", -- 0x11C8
    x"97",x"47",x"D6",x"4F",x"C1",x"80",x"22",x"11", -- 0x11D0
    x"8E",x"BD",x"C0",x"BD",x"BA",x"CA",x"96",x"47", -- 0x11D8
    x"80",x"09",x"20",x"EC",x"BD",x"BB",x"82",x"0C", -- 0x11E0
    x"47",x"8E",x"BD",x"BB",x"BD",x"BC",x"A0",x"2E", -- 0x11E8
    x"F3",x"8E",x"BD",x"B6",x"BD",x"BC",x"A0",x"2E", -- 0x11F0
    x"07",x"BD",x"BB",x"6A",x"0A",x"47",x"20",x"F1", -- 0x11F8
    x"35",x"C0",x"34",x"40",x"BD",x"B9",x"B4",x"BD", -- 0x1200
    x"BC",x"C8",x"35",x"40",x"8E",x"BE",x"C5",x"C6", -- 0x1208
    x"80",x"8D",x"36",x"96",x"53",x"AB",x"03",x"97", -- 0x1210
    x"53",x"96",x"52",x"A9",x"02",x"97",x"52",x"96", -- 0x1218
    x"51",x"A9",x"01",x"97",x"51",x"96",x"50",x"A9", -- 0x1220
    x"84",x"97",x"50",x"5C",x"56",x"59",x"28",x"E3", -- 0x1228
    x"24",x"03",x"C0",x"0B",x"50",x"CB",x"2F",x"30", -- 0x1230
    x"04",x"1F",x"98",x"84",x"7F",x"A7",x"C0",x"53", -- 0x1238
    x"C4",x"80",x"8C",x"BE",x"E9",x"26",x"CA",x"6F", -- 0x1240
    x"C4",x"0A",x"45",x"26",x"09",x"DF",x"39",x"86", -- 0x1248
    x"2E",x"A7",x"C0",x"0F",x"D7",x"39",x"0A",x"D7", -- 0x1250
    x"26",x"08",x"86",x"03",x"97",x"D7",x"86",x"2C", -- 0x1258
    x"A7",x"C0",x"39",x"96",x"47",x"8B",x"0A",x"97", -- 0x1260
    x"45",x"4C",x"80",x"03",x"24",x"FC",x"8B",x"05", -- 0x1268
    x"97",x"D7",x"96",x"DA",x"84",x"40",x"26",x"02", -- 0x1270
    x"97",x"D7",x"39",x"34",x"02",x"8D",x"CA",x"35", -- 0x1278
    x"02",x"4A",x"2B",x"0A",x"34",x"02",x"86",x"30", -- 0x1280
    x"A7",x"C0",x"A6",x"E0",x"26",x"ED",x"39",x"CE", -- 0x1288
    x"92",x"9C",x"96",x"B6",x"48",x"EE",x"C6",x"39", -- 0x1290
    x"8D",x"F5",x"6E",x"C4",x"92",x"A6",x"92",x"C2", -- 0x1298
    x"92",x"A6",x"92",x"C2",x"92",x"A6",x"34",x"44", -- 0x12A0
    x"D6",x"B9",x"96",x"C0",x"3D",x"D3",x"BA",x"1F", -- 0x12A8
    x"01",x"D6",x"BE",x"54",x"54",x"54",x"3A",x"96", -- 0x12B0
    x"BE",x"84",x"07",x"CE",x"92",x"DD",x"A6",x"C6", -- 0x12B8
    x"35",x"C4",x"34",x"44",x"D6",x"B9",x"96",x"C0", -- 0x12C0
    x"3D",x"D3",x"BA",x"1F",x"01",x"D6",x"BE",x"54", -- 0x12C8
    x"54",x"3A",x"96",x"BE",x"84",x"03",x"CE",x"92", -- 0x12D0
    x"E5",x"A6",x"C6",x"35",x"C4",x"80",x"40",x"20", -- 0x12D8
    x"10",x"08",x"04",x"02",x"01",x"C0",x"30",x"0C", -- 0x12E0
    x"03",x"D6",x"B9",x"3A",x"39",x"44",x"24",x"03", -- 0x12E8
    x"46",x"30",x"01",x"39",x"44",x"24",x"F6",x"86", -- 0x12F0
    x"C0",x"30",x"01",x"39",x"BD",x"B7",x"34",x"10", -- 0x12F8
    x"8E",x"00",x"BD",x"C1",x"C0",x"25",x"02",x"C6", -- 0x1300
    x"BF",x"4F",x"ED",x"22",x"DC",x"2B",x"10",x"83", -- 0x1308
    x"01",x"00",x"25",x"03",x"CC",x"00",x"FF",x"ED", -- 0x1310
    x"A4",x"39",x"BD",x"92",x"FC",x"CE",x"00",x"BD", -- 0x1318
    x"96",x"B6",x"81",x"02",x"24",x"06",x"EC",x"42", -- 0x1320
    x"44",x"56",x"ED",x"42",x"96",x"B6",x"81",x"04", -- 0x1328
    x"24",x"06",x"EC",x"C4",x"44",x"56",x"ED",x"C4", -- 0x1330
    x"39",x"BD",x"93",x"B2",x"BD",x"93",x"1D",x"BD", -- 0x1338
    x"92",x"98",x"A4",x"84",x"D6",x"B6",x"56",x"24", -- 0x1340
    x"12",x"81",x"04",x"25",x"04",x"46",x"46",x"20", -- 0x1348
    x"F8",x"4C",x"48",x"9B",x"C1",x"44",x"1F",x"89", -- 0x1350
    x"7E",x"B4",x"F3",x"4D",x"27",x"F8",x"4F",x"20", -- 0x1358
    x"F0",x"86",x"01",x"20",x"01",x"4F",x"97",x"C2", -- 0x1360
    x"BD",x"B2",x"6A",x"BD",x"93",x"1A",x"BD",x"95", -- 0x1368
    x"81",x"BD",x"B2",x"67",x"BD",x"92",x"98",x"E6", -- 0x1370
    x"84",x"34",x"04",x"1F",x"89",x"43",x"A4",x"84", -- 0x1378
    x"D4",x"B5",x"34",x"04",x"AA",x"E0",x"A7",x"84", -- 0x1380
    x"A0",x"E0",x"9A",x"DB",x"97",x"DB",x"39",x"9E", -- 0x1388
    x"C7",x"9F",x"BD",x"9E",x"C9",x"9F",x"BF",x"81", -- 0x1390
    x"AC",x"27",x"03",x"BD",x"93",x"B2",x"C6",x"AC", -- 0x1398
    x"BD",x"B2",x"6F",x"BD",x"B2",x"6A",x"BD",x"B7", -- 0x13A0
    x"34",x"10",x"8E",x"00",x"C3",x"BD",x"93",x"03", -- 0x13A8
    x"20",x"06",x"BD",x"B2",x"6A",x"BD",x"92",x"FC", -- 0x13B0
    x"7E",x"B2",x"67",x"81",x"89",x"10",x"27",x"F5", -- 0x13B8
    x"FF",x"81",x"28",x"27",x"09",x"81",x"AC",x"27", -- 0x13C0
    x"05",x"C6",x"40",x"BD",x"B2",x"6F",x"BD",x"93", -- 0x13C8
    x"8F",x"9E",x"C3",x"9F",x"C7",x"9E",x"C5",x"9F", -- 0x13D0
    x"C9",x"BD",x"B2",x"6D",x"81",x"BE",x"27",x"09", -- 0x13D8
    x"81",x"BD",x"10",x"26",x"1E",x"91",x"C6",x"01", -- 0x13E0
    x"86",x"5F",x"34",x"04",x"9D",x"9F",x"BD",x"94", -- 0x13E8
    x"20",x"35",x"04",x"D7",x"C2",x"BD",x"95",x"9A", -- 0x13F0
    x"9D",x"A5",x"10",x"27",x"00",x"A3",x"BD",x"B2", -- 0x13F8
    x"6D",x"C6",x"42",x"BD",x"B2",x"6F",x"26",x"21", -- 0x1400
    x"8D",x"3A",x"8D",x"62",x"9E",x"BD",x"34",x"10", -- 0x1408
    x"9E",x"C3",x"9F",x"BD",x"8D",x"58",x"35",x"10", -- 0x1410
    x"9F",x"BD",x"9E",x"C5",x"9F",x"BF",x"20",x"24", -- 0x1418
    x"BD",x"93",x"1D",x"CE",x"00",x"C3",x"7E",x"93", -- 0x1420
    x"20",x"C6",x"46",x"BD",x"B2",x"6F",x"20",x"04", -- 0x1428
    x"30",x"1F",x"9F",x"BF",x"BD",x"94",x"44",x"9E", -- 0x1430
    x"BF",x"9C",x"C5",x"27",x"06",x"24",x"F1",x"30", -- 0x1438
    x"01",x"20",x"EF",x"39",x"9E",x"BD",x"34",x"10", -- 0x1440
    x"BD",x"97",x"1D",x"24",x"04",x"9E",x"C3",x"9F", -- 0x1448
    x"BD",x"1F",x"02",x"31",x"21",x"BD",x"92",x"98", -- 0x1450
    x"35",x"40",x"DF",x"BD",x"8D",x"36",x"97",x"D7", -- 0x1458
    x"BD",x"93",x"77",x"96",x"D7",x"AD",x"C4",x"31", -- 0x1460
    x"3F",x"26",x"F3",x"39",x"35",x"06",x"DC",x"BF", -- 0x1468
    x"34",x"06",x"BD",x"97",x"10",x"24",x"04",x"9E", -- 0x1470
    x"C5",x"9F",x"BF",x"1F",x"02",x"31",x"21",x"BD", -- 0x1478
    x"92",x"98",x"35",x"40",x"DF",x"BF",x"8D",x"15", -- 0x1480
    x"20",x"D4",x"92",x"ED",x"92",x"F4",x"92",x"ED", -- 0x1488
    x"92",x"F4",x"92",x"ED",x"CE",x"94",x"8A",x"D6", -- 0x1490
    x"B6",x"58",x"EE",x"C5",x"39",x"CE",x"92",x"E9", -- 0x1498
    x"39",x"10",x"8E",x"95",x"0D",x"BD",x"97",x"10", -- 0x14A0
    x"10",x"27",x"FF",x"98",x"24",x"04",x"10",x"8E", -- 0x14A8
    x"95",x"1B",x"34",x"06",x"CE",x"95",x"06",x"BD", -- 0x14B0
    x"97",x"1D",x"27",x"B0",x"24",x"03",x"CE",x"95", -- 0x14B8
    x"14",x"10",x"A3",x"E4",x"35",x"10",x"24",x"04", -- 0x14C0
    x"1E",x"32",x"1E",x"01",x"34",x"46",x"34",x"06", -- 0x14C8
    x"44",x"56",x"25",x"09",x"11",x"83",x"95",x"0E", -- 0x14D0
    x"25",x"03",x"83",x"00",x"01",x"34",x"16",x"BD", -- 0x14D8
    x"92",x"8F",x"AD",x"C4",x"BD",x"93",x"77",x"AE", -- 0x14E0
    x"66",x"27",x"17",x"30",x"1F",x"AF",x"66",x"AD", -- 0x14E8
    x"F8",x"08",x"EC",x"E4",x"E3",x"62",x"ED",x"E4", -- 0x14F0
    x"A3",x"64",x"25",x"E6",x"ED",x"E4",x"AD",x"A4", -- 0x14F8
    x"20",x"E0",x"35",x"10",x"35",x"F6",x"9E",x"BD", -- 0x1500
    x"30",x"01",x"9F",x"BD",x"39",x"9E",x"BF",x"30", -- 0x1508
    x"01",x"9F",x"BF",x"39",x"9E",x"BD",x"30",x"1F", -- 0x1510
    x"9F",x"BD",x"39",x"9E",x"BF",x"30",x"1F",x"9F", -- 0x1518
    x"BF",x"39",x"CE",x"00",x"D3",x"8E",x"00",x"FF", -- 0x1520
    x"AF",x"C4",x"8E",x"00",x"BF",x"AF",x"42",x"7E", -- 0x1528
    x"93",x"20",x"27",x"0E",x"8D",x"24",x"86",x"55", -- 0x1530
    x"3D",x"9E",x"BA",x"E7",x"80",x"9C",x"B7",x"26", -- 0x1538
    x"FA",x"39",x"D6",x"B3",x"20",x"F0",x"81",x"2C", -- 0x1540
    x"27",x"08",x"8D",x"0E",x"D7",x"B2",x"9D",x"A5", -- 0x1548
    x"27",x"07",x"BD",x"B2",x"6D",x"8D",x"03",x"D7", -- 0x1550
    x"B3",x"39",x"BD",x"B7",x"0B",x"C1",x"09",x"10", -- 0x1558
    x"24",x"1E",x"E7",x"4F",x"C1",x"05",x"25",x"04", -- 0x1560
    x"86",x"08",x"C0",x"04",x"34",x"02",x"96",x"B6", -- 0x1568
    x"46",x"24",x"08",x"5D",x"26",x"02",x"C6",x"04", -- 0x1570
    x"5A",x"35",x"82",x"56",x"25",x"F8",x"5F",x"20", -- 0x1578
    x"F8",x"BD",x"95",x"9A",x"9D",x"A5",x"27",x"10", -- 0x1580
    x"81",x"29",x"27",x"0C",x"BD",x"B2",x"6D",x"81", -- 0x1588
    x"2C",x"27",x"05",x"BD",x"95",x"5A",x"8D",x"0A", -- 0x1590
    x"0E",x"A5",x"D6",x"B2",x"0D",x"C2",x"26",x"02", -- 0x1598
    x"D6",x"B3",x"D7",x"B4",x"86",x"55",x"3D",x"D7", -- 0x15A0
    x"B5",x"39",x"26",x"23",x"34",x"16",x"8E",x"FF", -- 0x15A8
    x"C8",x"A7",x"0A",x"A7",x"08",x"A7",x"06",x"A7", -- 0x15B0
    x"04",x"A7",x"02",x"A7",x"01",x"A7",x"1E",x"A7", -- 0x15B8
    x"1C",x"A7",x"1A",x"A7",x"18",x"B6",x"FF",x"22", -- 0x15C0
    x"84",x"07",x"B7",x"FF",x"22",x"35",x"96",x"34", -- 0x15C8
    x"16",x"96",x"B6",x"8B",x"03",x"C6",x"10",x"3D", -- 0x15D0
    x"CA",x"80",x"DA",x"C1",x"B6",x"FF",x"22",x"84", -- 0x15D8
    x"07",x"34",x"02",x"EA",x"E0",x"F7",x"FF",x"22", -- 0x15E0
    x"96",x"BA",x"44",x"BD",x"96",x"0F",x"96",x"B6", -- 0x15E8
    x"8B",x"03",x"81",x"07",x"26",x"01",x"4A",x"8D", -- 0x15F0
    x"02",x"35",x"96",x"C6",x"03",x"8E",x"FF",x"C0", -- 0x15F8
    x"46",x"24",x"04",x"A7",x"01",x"20",x"02",x"A7", -- 0x1600
    x"84",x"30",x"02",x"5A",x"26",x"F2",x"39",x"C6", -- 0x1608
    x"07",x"8E",x"FF",x"C6",x"20",x"EA",x"B6",x"FF", -- 0x1610
    x"22",x"84",x"F7",x"9A",x"C1",x"B7",x"FF",x"22", -- 0x1618
    x"39",x"81",x"2C",x"27",x"2B",x"BD",x"B7",x"0B", -- 0x1620
    x"C1",x"05",x"24",x"41",x"96",x"BC",x"97",x"BA", -- 0x1628
    x"58",x"CE",x"97",x"07",x"AB",x"C5",x"91",x"19", -- 0x1630
    x"22",x"33",x"97",x"B7",x"33",x"5F",x"A6",x"C5", -- 0x1638
    x"97",x"B9",x"54",x"D7",x"B6",x"4F",x"97",x"B3", -- 0x1640
    x"86",x"03",x"97",x"B2",x"9D",x"A5",x"27",x"1C", -- 0x1648
    x"BD",x"B7",x"38",x"5D",x"27",x"17",x"5A",x"86", -- 0x1650
    x"06",x"3D",x"DB",x"BC",x"34",x"04",x"DB",x"B7", -- 0x1658
    x"D0",x"BA",x"D1",x"19",x"22",x"07",x"D7",x"B7", -- 0x1660
    x"35",x"04",x"D7",x"BA",x"39",x"7E",x"B4",x"4A", -- 0x1668
    x"81",x"2C",x"27",x"0B",x"BD",x"B7",x"0B",x"5D", -- 0x1670
    x"BD",x"95",x"AA",x"9D",x"A5",x"27",x"ED",x"BD", -- 0x1678
    x"B7",x"38",x"5D",x"27",x"02",x"C6",x"08",x"D7", -- 0x1680
    x"C1",x"20",x"8B",x"BD",x"B7",x"0B",x"5D",x"27", -- 0x1688
    x"DC",x"C1",x"09",x"24",x"D8",x"86",x"06",x"3D", -- 0x1690
    x"DB",x"BC",x"1F",x"98",x"C6",x"01",x"1F",x"02", -- 0x1698
    x"10",x"93",x"B7",x"25",x"C8",x"93",x"19",x"D3", -- 0x16A0
    x"1B",x"1F",x"01",x"4C",x"93",x"21",x"24",x"BD", -- 0x16A8
    x"BD",x"80",x"D0",x"12",x"DE",x"1B",x"9F",x"1B", -- 0x16B0
    x"11",x"93",x"1B",x"24",x"17",x"A6",x"C2",x"A7", -- 0x16B8
    x"82",x"11",x"93",x"19",x"26",x"F7",x"10",x"9F", -- 0x16C0
    x"19",x"6F",x"3F",x"BD",x"AC",x"EF",x"BD",x"AD", -- 0x16C8
    x"26",x"7E",x"AD",x"9E",x"DE",x"19",x"10",x"9F", -- 0x16D0
    x"19",x"6F",x"3F",x"A6",x"C0",x"A7",x"A0",x"10", -- 0x16D8
    x"9C",x"1B",x"26",x"F7",x"20",x"E5",x"C6",x"1E", -- 0x16E0
    x"D7",x"19",x"86",x"06",x"97",x"BC",x"97",x"BA", -- 0x16E8
    x"4F",x"97",x"B6",x"86",x"10",x"97",x"B9",x"86", -- 0x16F0
    x"03",x"97",x"B2",x"86",x"0C",x"97",x"B7",x"9E", -- 0x16F8
    x"19",x"6F",x"1F",x"7E",x"AD",x"19",x"10",x"06", -- 0x1700
    x"20",x"0C",x"10",x"0C",x"20",x"18",x"20",x"18", -- 0x1708
    x"DC",x"C5",x"93",x"BF",x"24",x"3B",x"34",x"01", -- 0x1710
    x"BD",x"9D",x"C3",x"35",x"81",x"DC",x"C3",x"93", -- 0x1718
    x"BD",x"20",x"F1",x"8D",x"1A",x"34",x"06",x"C6", -- 0x1720
    x"A5",x"BD",x"B2",x"6F",x"8D",x"11",x"35",x"10", -- 0x1728
    x"1F",x"03",x"10",x"8E",x"03",x"00",x"EC",x"81", -- 0x1730
    x"ED",x"C1",x"31",x"3F",x"26",x"F8",x"39",x"BD", -- 0x1738
    x"B7",x"0B",x"5D",x"27",x"0D",x"D1",x"19",x"22", -- 0x1740
    x"09",x"5A",x"86",x"06",x"3D",x"DB",x"BC",x"1E", -- 0x1748
    x"89",x"39",x"7E",x"B4",x"4A",x"5F",x"20",x"02", -- 0x1750
    x"C6",x"01",x"D7",x"D8",x"BD",x"01",x"A0",x"81", -- 0x1758
    x"40",x"26",x"02",x"9D",x"9F",x"BD",x"93",x"8F", -- 0x1760
    x"BD",x"B2",x"6D",x"BD",x"98",x"CC",x"1F",x"10", -- 0x1768
    x"EE",x"84",x"33",x"5E",x"33",x"CB",x"DF",x"D1", -- 0x1770
    x"30",x"02",x"E6",x"84",x"58",x"3A",x"9F",x"CF", -- 0x1778
    x"96",x"06",x"26",x"CE",x"0F",x"D4",x"9D",x"A5", -- 0x1780
    x"27",x"2D",x"03",x"D4",x"BD",x"B2",x"6D",x"0D", -- 0x1788
    x"D8",x"26",x"07",x"C6",x"47",x"BD",x"B2",x"6F", -- 0x1790
    x"20",x"30",x"C6",x"05",x"8E",x"98",x"39",x"EE", -- 0x1798
    x"81",x"10",x"AE",x"81",x"A1",x"80",x"27",x"06", -- 0x17A0
    x"5A",x"26",x"F4",x"7E",x"B2",x"77",x"10",x"9F", -- 0x17A8
    x"D5",x"DF",x"D9",x"9D",x"9F",x"20",x"13",x"C6", -- 0x17B0
    x"F8",x"96",x"B6",x"46",x"24",x"02",x"C6",x"FC", -- 0x17B8
    x"1F",x"98",x"D4",x"BE",x"D7",x"BE",x"94",x"C4", -- 0x17C0
    x"97",x"C4",x"BD",x"97",x"1D",x"24",x"04",x"9E", -- 0x17C8
    x"C3",x"9F",x"BD",x"DD",x"C3",x"BD",x"97",x"10", -- 0x17D0
    x"24",x"04",x"9E",x"C5",x"9F",x"BF",x"DD",x"C5", -- 0x17D8
    x"96",x"B6",x"46",x"DC",x"C3",x"24",x"04",x"D3", -- 0x17E0
    x"C3",x"DD",x"C3",x"BD",x"94",x"20",x"DC",x"C3", -- 0x17E8
    x"9E",x"C5",x"30",x"01",x"9F",x"C5",x"0D",x"D4", -- 0x17F0
    x"26",x"58",x"44",x"56",x"44",x"56",x"44",x"56", -- 0x17F8
    x"C3",x"00",x"01",x"DD",x"C3",x"BD",x"92",x"98", -- 0x1800
    x"D6",x"C4",x"34",x"10",x"0D",x"D8",x"27",x"21", -- 0x1808
    x"8D",x"11",x"A6",x"C4",x"A7",x"80",x"5A",x"26", -- 0x1810
    x"F3",x"35",x"10",x"BD",x"92",x"E9",x"0A",x"C6", -- 0x1818
    x"26",x"E6",x"39",x"DE",x"CF",x"33",x"41",x"DF", -- 0x1820
    x"CF",x"11",x"93",x"D1",x"26",x"F4",x"7E",x"B4", -- 0x1828
    x"4A",x"A6",x"80",x"8D",x"EE",x"A7",x"C4",x"20", -- 0x1830
    x"DD",x"98",x"94",x"98",x"9B",x"BD",x"98",x"9B", -- 0x1838
    x"98",x"94",x"BE",x"98",x"B1",x"98",x"9B",x"B1", -- 0x1840
    x"98",x"94",x"98",x"B1",x"B0",x"98",x"A1",x"98", -- 0x1848
    x"A1",x"A8",x"C3",x"00",x"01",x"DD",x"C3",x"96", -- 0x1850
    x"D8",x"26",x"09",x"DE",x"D1",x"A7",x"C2",x"11", -- 0x1858
    x"93",x"CF",x"22",x"F9",x"BD",x"92",x"98",x"D6", -- 0x1860
    x"B6",x"56",x"24",x"02",x"84",x"AA",x"C6",x"01", -- 0x1868
    x"10",x"9E",x"CF",x"34",x"12",x"DE",x"C3",x"34", -- 0x1870
    x"42",x"54",x"24",x"08",x"56",x"31",x"21",x"10", -- 0x1878
    x"9C",x"D1",x"27",x"AA",x"0D",x"D8",x"27",x"1F", -- 0x1880
    x"E5",x"A4",x"27",x"04",x"6E",x"9F",x"00",x"D5", -- 0x1888
    x"6E",x"9F",x"00",x"D9",x"43",x"A4",x"84",x"A7", -- 0x1890
    x"84",x"20",x"16",x"AA",x"84",x"A7",x"84",x"20", -- 0x1898
    x"10",x"A8",x"84",x"A7",x"84",x"20",x"0A",x"A5", -- 0x18A0
    x"84",x"27",x"06",x"1F",x"98",x"AA",x"A4",x"A7", -- 0x18A8
    x"A4",x"35",x"42",x"BD",x"92",x"ED",x"33",x"5F", -- 0x18B0
    x"11",x"93",x"8A",x"26",x"BA",x"AE",x"61",x"96", -- 0x18B8
    x"B9",x"30",x"86",x"35",x"02",x"32",x"62",x"0A", -- 0x18C0
    x"C6",x"26",x"A8",x"39",x"BD",x"B3",x"57",x"E6", -- 0x18C8
    x"82",x"A6",x"82",x"1F",x"03",x"9E",x"1D",x"9C", -- 0x18D0
    x"1F",x"10",x"27",x"1B",x"6D",x"11",x"A3",x"84", -- 0x18D8
    x"27",x"06",x"EC",x"02",x"30",x"8B",x"20",x"EF", -- 0x18E0
    x"30",x"02",x"39",x"39",x"81",x"40",x"26",x"02", -- 0x18E8
    x"9D",x"9F",x"BD",x"93",x"B2",x"BD",x"93",x"1D", -- 0x18F0
    x"86",x"01",x"97",x"C2",x"BD",x"95",x"81",x"DC", -- 0x18F8
    x"B4",x"34",x"06",x"9D",x"A5",x"27",x"03",x"BD", -- 0x1900
    x"95",x"81",x"96",x"B5",x"97",x"D8",x"35",x"06", -- 0x1908
    x"DD",x"B4",x"4F",x"34",x"56",x"BD",x"95",x"22", -- 0x1910
    x"BD",x"92",x"8F",x"DF",x"D9",x"BD",x"99",x"DF", -- 0x1918
    x"27",x"0F",x"BD",x"99",x"CB",x"86",x"01",x"97", -- 0x1920
    x"D7",x"BD",x"99",x"BA",x"00",x"D7",x"BD",x"99", -- 0x1928
    x"BA",x"10",x"DF",x"DC",x"0D",x"DB",x"26",x"03", -- 0x1930
    x"10",x"DE",x"DC",x"35",x"56",x"0F",x"DB",x"10", -- 0x1938
    x"DF",x"DC",x"30",x"01",x"9F",x"BD",x"DF",x"D1", -- 0x1940
    x"97",x"D7",x"27",x"9F",x"2B",x"06",x"5C",x"D1", -- 0x1948
    x"D6",x"23",x"05",x"5F",x"5D",x"27",x"DD",x"5A", -- 0x1950
    x"D7",x"C0",x"BD",x"99",x"DF",x"27",x"0F",x"10", -- 0x1958
    x"83",x"00",x"03",x"25",x"04",x"30",x"1E",x"8D", -- 0x1960
    x"38",x"BD",x"99",x"CB",x"8D",x"4C",x"43",x"53", -- 0x1968
    x"D3",x"D1",x"DD",x"D1",x"2F",x"16",x"BD",x"95", -- 0x1970
    x"06",x"BD",x"9A",x"12",x"26",x"05",x"CC",x"FF", -- 0x1978
    x"FF",x"20",x"ED",x"BD",x"95",x"14",x"8D",x"3E", -- 0x1980
    x"8D",x"5E",x"20",x"E0",x"BD",x"95",x"06",x"30", -- 0x1988
    x"8B",x"9F",x"BD",x"43",x"53",x"83",x"00",x"01", -- 0x1990
    x"2F",x"04",x"1F",x"01",x"8D",x"03",x"7E",x"99", -- 0x1998
    x"34",x"DD",x"CB",x"35",x"20",x"DC",x"BD",x"34", -- 0x19A0
    x"16",x"96",x"D7",x"40",x"D6",x"C0",x"34",x"06", -- 0x19A8
    x"34",x"20",x"C6",x"02",x"BD",x"AC",x"33",x"DC", -- 0x19B0
    x"CB",x"39",x"DD",x"CB",x"35",x"20",x"DC",x"C3", -- 0x19B8
    x"34",x"16",x"96",x"D7",x"20",x"E6",x"9E",x"BD", -- 0x19C0
    x"9F",x"C3",x"39",x"DD",x"CD",x"10",x"9E",x"C3", -- 0x19C8
    x"8D",x"F4",x"10",x"9F",x"BD",x"8D",x"11",x"9E", -- 0x19D0
    x"CD",x"30",x"8B",x"C3",x"00",x"01",x"39",x"BD", -- 0x19D8
    x"99",x"C6",x"10",x"8E",x"95",x"14",x"20",x"06", -- 0x19E0
    x"10",x"8E",x"95",x"06",x"AD",x"A4",x"DE",x"8A", -- 0x19E8
    x"9E",x"BD",x"2B",x"17",x"9C",x"D3",x"22",x"13", -- 0x19F0
    x"34",x"60",x"8D",x"16",x"27",x"0B",x"BD",x"93", -- 0x19F8
    x"77",x"35",x"60",x"33",x"41",x"AD",x"A4",x"20", -- 0x1A00
    x"E9",x"35",x"60",x"1F",x"30",x"1F",x"01",x"93", -- 0x1A08
    x"8A",x"39",x"AD",x"9F",x"00",x"D9",x"1F",x"89", -- 0x1A10
    x"D4",x"D8",x"34",x"06",x"A4",x"84",x"A1",x"61", -- 0x1A18
    x"35",x"86",x"9E",x"8A",x"C6",x"01",x"34",x"14", -- 0x1A20
    x"BD",x"B1",x"56",x"5F",x"BD",x"A9",x"A2",x"BD", -- 0x1A28
    x"A9",x"76",x"BD",x"B6",x"54",x"20",x"02",x"35", -- 0x1A30
    x"14",x"D7",x"D8",x"27",x"FA",x"9F",x"D9",x"10", -- 0x1A38
    x"27",x"0F",x"31",x"0D",x"D8",x"27",x"F0",x"BD", -- 0x1A40
    x"9B",x"98",x"81",x"3B",x"27",x"F5",x"81",x"27", -- 0x1A48
    x"27",x"F1",x"81",x"58",x"10",x"27",x"01",x"B2", -- 0x1A50
    x"8D",x"02",x"20",x"E7",x"81",x"4F",x"26",x"0D", -- 0x1A58
    x"D6",x"DE",x"5C",x"8D",x"5B",x"5A",x"C1",x"04", -- 0x1A60
    x"22",x"63",x"D7",x"DE",x"39",x"81",x"56",x"26", -- 0x1A68
    x"1A",x"D6",x"DF",x"54",x"54",x"C0",x"1F",x"8D", -- 0x1A70
    x"47",x"C1",x"1F",x"22",x"50",x"58",x"58",x"34", -- 0x1A78
    x"04",x"CC",x"7E",x"7E",x"AB",x"E4",x"E0",x"E0", -- 0x1A80
    x"DD",x"DF",x"39",x"81",x"4C",x"26",x"23",x"D6", -- 0x1A88
    x"E1",x"8D",x"2D",x"5D",x"27",x"37",x"D7",x"E1", -- 0x1A90
    x"0F",x"E5",x"8D",x"03",x"24",x"FC",x"39",x"0D", -- 0x1A98
    x"D8",x"27",x"0A",x"BD",x"9B",x"98",x"81",x"2E", -- 0x1AA0
    x"27",x"05",x"BD",x"9B",x"E2",x"43",x"39",x"0C", -- 0x1AA8
    x"E5",x"39",x"81",x"54",x"26",x"0D",x"D6",x"E2", -- 0x1AB0
    x"8D",x"06",x"5D",x"27",x"10",x"D7",x"E2",x"39", -- 0x1AB8
    x"7E",x"9B",x"AC",x"81",x"50",x"26",x"24",x"BD", -- 0x1AC0
    x"9C",x"CB",x"5D",x"26",x"03",x"7E",x"B4",x"4A", -- 0x1AC8
    x"96",x"E5",x"9E",x"DF",x"34",x"12",x"86",x"7E", -- 0x1AD0
    x"97",x"DF",x"97",x"E0",x"0F",x"E5",x"8D",x"07", -- 0x1AD8
    x"35",x"12",x"97",x"E5",x"9F",x"DF",x"39",x"6F", -- 0x1AE0
    x"E2",x"20",x"40",x"81",x"4E",x"26",x"03",x"BD", -- 0x1AE8
    x"9B",x"98",x"81",x"41",x"25",x"04",x"81",x"47", -- 0x1AF0
    x"23",x"05",x"BD",x"9B",x"BE",x"20",x"23",x"80", -- 0x1AF8
    x"41",x"8E",x"9C",x"5B",x"E6",x"86",x"0D",x"D8", -- 0x1B00
    x"27",x"18",x"BD",x"9B",x"98",x"81",x"23",x"27", -- 0x1B08
    x"04",x"81",x"2B",x"26",x"03",x"5C",x"20",x"0A", -- 0x1B10
    x"81",x"2D",x"26",x"03",x"5A",x"20",x"03",x"BD", -- 0x1B18
    x"9B",x"E2",x"5A",x"C1",x"0B",x"22",x"A6",x"34", -- 0x1B20
    x"04",x"D6",x"E1",x"96",x"E2",x"3D",x"DD",x"D5", -- 0x1B28
    x"33",x"61",x"96",x"DE",x"81",x"01",x"22",x"2C", -- 0x1B30
    x"8E",x"9C",x"62",x"C6",x"18",x"3D",x"3A",x"35", -- 0x1B38
    x"04",x"58",x"3A",x"31",x"84",x"8D",x"45",x"DD", -- 0x1B40
    x"E3",x"8D",x"0C",x"96",x"DF",x"8D",x"0B",x"8D", -- 0x1B48
    x"06",x"96",x"E0",x"8D",x"05",x"20",x"F2",x"86", -- 0x1B50
    x"7E",x"12",x"B7",x"FF",x"20",x"AE",x"A4",x"30", -- 0x1B58
    x"1F",x"26",x"FC",x"39",x"8E",x"9C",x"7A",x"C6", -- 0x1B60
    x"0C",x"3D",x"3A",x"35",x"04",x"3A",x"8D",x"1C", -- 0x1B68
    x"DD",x"E3",x"8D",x"0C",x"96",x"DF",x"8D",x"0B", -- 0x1B70
    x"8D",x"06",x"96",x"E0",x"8D",x"05",x"20",x"F2", -- 0x1B78
    x"86",x"7E",x"12",x"B7",x"FF",x"20",x"A6",x"84", -- 0x1B80
    x"4A",x"26",x"FD",x"39",x"C6",x"FF",x"96",x"E5", -- 0x1B88
    x"27",x"05",x"8B",x"02",x"3D",x"44",x"56",x"39", -- 0x1B90
    x"34",x"10",x"0D",x"D8",x"27",x"4D",x"9E",x"D9", -- 0x1B98
    x"A6",x"80",x"9F",x"D9",x"0A",x"D8",x"81",x"20", -- 0x1BA0
    x"27",x"F0",x"35",x"90",x"8D",x"EA",x"81",x"2B", -- 0x1BA8
    x"27",x"3C",x"81",x"2D",x"27",x"3C",x"81",x"3E", -- 0x1BB0
    x"27",x"42",x"81",x"3C",x"27",x"39",x"81",x"3D", -- 0x1BB8
    x"27",x"3F",x"BD",x"90",x"AA",x"25",x"24",x"5F", -- 0x1BC0
    x"80",x"30",x"97",x"D7",x"86",x"0A",x"3D",x"4D", -- 0x1BC8
    x"26",x"19",x"DB",x"D7",x"25",x"15",x"0D",x"D8", -- 0x1BD0
    x"27",x"17",x"BD",x"9B",x"98",x"BD",x"90",x"AA", -- 0x1BD8
    x"24",x"E6",x"0C",x"D8",x"9E",x"D9",x"30",x"1F", -- 0x1BE0
    x"9F",x"D9",x"39",x"7E",x"B4",x"4A",x"5C",x"27", -- 0x1BE8
    x"FA",x"39",x"5D",x"27",x"F6",x"5A",x"39",x"5D", -- 0x1BF0
    x"27",x"F1",x"54",x"39",x"5D",x"2B",x"EC",x"58", -- 0x1BF8
    x"39",x"34",x"60",x"8D",x"16",x"BD",x"B7",x"0E", -- 0x1C00
    x"35",x"E0",x"BD",x"9C",x"1B",x"C6",x"02",x"BD", -- 0x1C08
    x"AC",x"33",x"D6",x"D8",x"9E",x"D9",x"34",x"14", -- 0x1C10
    x"7E",x"9A",x"32",x"9E",x"D9",x"34",x"10",x"BD", -- 0x1C18
    x"9B",x"98",x"BD",x"B3",x"A2",x"25",x"C4",x"BD", -- 0x1C20
    x"9B",x"98",x"81",x"3B",x"26",x"F9",x"35",x"10", -- 0x1C28
    x"DE",x"A6",x"34",x"40",x"9F",x"A6",x"BD",x"B2", -- 0x1C30
    x"84",x"35",x"10",x"9F",x"A6",x"39",x"4F",x"1F", -- 0x1C38
    x"8B",x"DC",x"E3",x"10",x"27",x"0D",x"74",x"93", -- 0x1C40
    x"D5",x"DD",x"E3",x"22",x"0D",x"0F",x"E3",x"0F", -- 0x1C48
    x"E4",x"35",x"02",x"10",x"EE",x"67",x"84",x"7F", -- 0x1C50
    x"34",x"02",x"3B",x"0A",x"0C",x"01",x"03",x"05", -- 0x1C58
    x"06",x"08",x"01",x"A8",x"01",x"90",x"01",x"7A", -- 0x1C60
    x"01",x"64",x"01",x"50",x"01",x"3D",x"01",x"2B", -- 0x1C68
    x"01",x"1A",x"01",x"0A",x"00",x"FB",x"00",x"ED", -- 0x1C70
    x"00",x"DF",x"00",x"D3",x"00",x"C7",x"00",x"BB", -- 0x1C78
    x"00",x"B1",x"00",x"A6",x"00",x"9D",x"00",x"94", -- 0x1C80
    x"00",x"8B",x"00",x"83",x"00",x"7C",x"00",x"75", -- 0x1C88
    x"00",x"6E",x"A6",x"9C",x"93",x"8B",x"83",x"7B", -- 0x1C90
    x"74",x"6D",x"67",x"61",x"5B",x"56",x"51",x"4C", -- 0x1C98
    x"47",x"43",x"3F",x"3B",x"37",x"34",x"31",x"2E", -- 0x1CA0
    x"2B",x"28",x"26",x"23",x"21",x"1F",x"1D",x"1B", -- 0x1CA8
    x"19",x"18",x"16",x"14",x"13",x"12",x"9E",x"8A", -- 0x1CB0
    x"C6",x"01",x"34",x"14",x"D7",x"C2",x"9F",x"D5", -- 0x1CB8
    x"BD",x"95",x"9A",x"BD",x"B1",x"56",x"BD",x"B6", -- 0x1CC0
    x"54",x"20",x"08",x"BD",x"9B",x"98",x"7E",x"9B", -- 0x1CC8
    x"BE",x"35",x"14",x"D7",x"D8",x"27",x"FA",x"9F", -- 0x1CD0
    x"D9",x"10",x"27",x"00",x"EA",x"0D",x"D8",x"27", -- 0x1CD8
    x"F0",x"BD",x"9B",x"98",x"81",x"3B",x"27",x"F5", -- 0x1CE0
    x"81",x"27",x"27",x"F1",x"81",x"4E",x"26",x"04", -- 0x1CE8
    x"03",x"D5",x"20",x"E9",x"81",x"42",x"26",x"04", -- 0x1CF0
    x"03",x"D6",x"20",x"E1",x"81",x"58",x"10",x"27", -- 0x1CF8
    x"00",x"96",x"81",x"4D",x"10",x"27",x"01",x"2A", -- 0x1D00
    x"34",x"02",x"C6",x"01",x"0D",x"D8",x"27",x"11", -- 0x1D08
    x"BD",x"9B",x"98",x"BD",x"B3",x"A2",x"34",x"01", -- 0x1D10
    x"BD",x"9B",x"E2",x"35",x"01",x"24",x"02",x"8D", -- 0x1D18
    x"AA",x"35",x"02",x"81",x"43",x"27",x"28",x"81", -- 0x1D20
    x"41",x"27",x"2E",x"81",x"53",x"27",x"32",x"81", -- 0x1D28
    x"55",x"27",x"5C",x"81",x"44",x"27",x"55",x"81", -- 0x1D30
    x"4C",x"27",x"4C",x"81",x"52",x"27",x"43",x"80", -- 0x1D38
    x"45",x"27",x"2F",x"4A",x"27",x"27",x"4A",x"27", -- 0x1D40
    x"32",x"4A",x"27",x"1D",x"7E",x"B4",x"4A",x"BD", -- 0x1D48
    x"95",x"5D",x"D7",x"B2",x"BD",x"95",x"9A",x"20", -- 0x1D50
    x"84",x"C1",x"04",x"24",x"EF",x"D7",x"E8",x"20", -- 0x1D58
    x"F6",x"C1",x"3F",x"24",x"E7",x"D7",x"E9",x"20", -- 0x1D60
    x"EE",x"4F",x"8D",x"58",x"21",x"4F",x"1F",x"01", -- 0x1D68
    x"20",x"59",x"4F",x"1F",x"01",x"8D",x"4D",x"1E", -- 0x1D70
    x"01",x"20",x"50",x"4F",x"1F",x"01",x"8D",x"44", -- 0x1D78
    x"20",x"49",x"4F",x"9E",x"8A",x"20",x"44",x"4F", -- 0x1D80
    x"8D",x"3A",x"20",x"F7",x"4F",x"20",x"03",x"4F", -- 0x1D88
    x"8D",x"32",x"9E",x"8A",x"1E",x"10",x"20",x"33", -- 0x1D90
    x"BD",x"9C",x"1B",x"C6",x"02",x"BD",x"AC",x"33", -- 0x1D98
    x"D6",x"D8",x"9E",x"D9",x"34",x"14",x"7E",x"9C", -- 0x1DA0
    x"C6",x"D6",x"E9",x"27",x"1B",x"4F",x"1E",x"01", -- 0x1DA8
    x"A7",x"E2",x"2A",x"02",x"8D",x"0D",x"BD",x"9F", -- 0x1DB0
    x"B5",x"1F",x"30",x"44",x"56",x"44",x"56",x"6D", -- 0x1DB8
    x"E0",x"2A",x"04",x"40",x"50",x"82",x"00",x"39", -- 0x1DC0
    x"1F",x"10",x"39",x"34",x"06",x"8D",x"DA",x"35", -- 0x1DC8
    x"10",x"34",x"06",x"8D",x"D4",x"35",x"10",x"10", -- 0x1DD0
    x"9E",x"E8",x"34",x"20",x"6D",x"E4",x"27",x"08", -- 0x1DD8
    x"1E",x"10",x"8D",x"DF",x"6A",x"E4",x"20",x"F4", -- 0x1DE0
    x"35",x"20",x"DE",x"8A",x"D3",x"C7",x"2B",x"02", -- 0x1DE8
    x"1F",x"03",x"1F",x"10",x"9E",x"8A",x"D3",x"C9", -- 0x1DF0
    x"2B",x"02",x"1F",x"01",x"11",x"83",x"01",x"00", -- 0x1DF8
    x"25",x"03",x"CE",x"00",x"FF",x"8C",x"00",x"C0", -- 0x1E00
    x"25",x"03",x"8E",x"00",x"BF",x"DC",x"C7",x"DD", -- 0x1E08
    x"BD",x"DC",x"C9",x"DD",x"BF",x"9F",x"C5",x"DF", -- 0x1E10
    x"C3",x"0D",x"D5",x"26",x"04",x"9F",x"C9",x"DF", -- 0x1E18
    x"C7",x"BD",x"94",x"20",x"0D",x"D6",x"26",x"03", -- 0x1E20
    x"BD",x"94",x"A1",x"0F",x"D5",x"0F",x"D6",x"7E", -- 0x1E28
    x"9C",x"DD",x"BD",x"9B",x"98",x"34",x"02",x"BD", -- 0x1E30
    x"9E",x"5E",x"34",x"06",x"BD",x"9B",x"98",x"81", -- 0x1E38
    x"2C",x"10",x"26",x"FF",x"07",x"BD",x"9E",x"5B", -- 0x1E40
    x"1F",x"01",x"35",x"40",x"35",x"02",x"81",x"2B", -- 0x1E48
    x"27",x"04",x"81",x"2D",x"26",x"A6",x"1F",x"30", -- 0x1E50
    x"7E",x"9D",x"CB",x"BD",x"9B",x"98",x"81",x"2B", -- 0x1E58
    x"27",x"07",x"81",x"2D",x"27",x"04",x"BD",x"9B", -- 0x1E60
    x"E2",x"4F",x"34",x"02",x"BD",x"9C",x"CB",x"35", -- 0x1E68
    x"02",x"4D",x"27",x"04",x"4F",x"50",x"82",x"00", -- 0x1E70
    x"39",x"00",x"00",x"00",x"01",x"FE",x"C5",x"19", -- 0x1E78
    x"19",x"FB",x"16",x"31",x"F2",x"F4",x"FB",x"4A", -- 0x1E80
    x"51",x"EC",x"84",x"61",x"F9",x"E1",x"C7",x"78", -- 0x1E88
    x"AE",x"D4",x"DC",x"8E",x"3B",x"C5",x"E5",x"A2", -- 0x1E90
    x"69",x"B5",x"06",x"B5",x"06",x"81",x"40",x"26", -- 0x1E98
    x"02",x"9D",x"9F",x"BD",x"95",x"22",x"BD",x"93", -- 0x1EA0
    x"B2",x"BD",x"93",x"1D",x"AE",x"C4",x"9F",x"CB", -- 0x1EA8
    x"AE",x"42",x"9F",x"CD",x"BD",x"B2",x"6D",x"BD", -- 0x1EB0
    x"B7",x"3D",x"CE",x"00",x"CF",x"AF",x"C4",x"BD", -- 0x1EB8
    x"93",x"20",x"86",x"01",x"97",x"C2",x"BD",x"95", -- 0x1EC0
    x"81",x"8E",x"01",x"00",x"9D",x"A5",x"27",x"0F", -- 0x1EC8
    x"BD",x"B2",x"6D",x"BD",x"B1",x"41",x"96",x"4F", -- 0x1ED0
    x"8B",x"08",x"97",x"4F",x"BD",x"B7",x"40",x"96", -- 0x1ED8
    x"B6",x"85",x"02",x"27",x"04",x"1F",x"10",x"30", -- 0x1EE0
    x"8B",x"9F",x"D1",x"C6",x"01",x"D7",x"C2",x"D7", -- 0x1EE8
    x"D8",x"BD",x"9F",x"E2",x"34",x"06",x"BD",x"9F", -- 0x1EF0
    x"E2",x"DD",x"D9",x"35",x"06",x"34",x"06",x"9E", -- 0x1EF8
    x"C3",x"9F",x"BD",x"9E",x"C5",x"9F",x"BF",x"CE", -- 0x1F00
    x"9E",x"7B",x"84",x"01",x"27",x"03",x"50",x"CB", -- 0x1F08
    x"08",x"58",x"58",x"33",x"C5",x"34",x"40",x"BD", -- 0x1F10
    x"9F",x"A7",x"35",x"40",x"33",x"5E",x"34",x"10", -- 0x1F18
    x"BD",x"9F",x"A7",x"35",x"20",x"A6",x"E4",x"84", -- 0x1F20
    x"03",x"27",x"06",x"81",x"03",x"27",x"02",x"1E", -- 0x1F28
    x"12",x"9F",x"C3",x"1F",x"21",x"DC",x"D1",x"BD", -- 0x1F30
    x"9F",x"B5",x"1F",x"20",x"4D",x"10",x"26",x"15", -- 0x1F38
    x"09",x"D7",x"C5",x"1F",x"30",x"97",x"C6",x"A6", -- 0x1F40
    x"E4",x"81",x"02",x"25",x"0E",x"81",x"06",x"24", -- 0x1F48
    x"0A",x"DC",x"CB",x"93",x"C3",x"24",x"11",x"4F", -- 0x1F50
    x"5F",x"20",x"0D",x"DC",x"CB",x"D3",x"C3",x"25", -- 0x1F58
    x"05",x"10",x"93",x"D3",x"25",x"02",x"DC",x"D3", -- 0x1F60
    x"DD",x"C3",x"A6",x"E4",x"81",x"04",x"25",x"0A", -- 0x1F68
    x"DC",x"CD",x"93",x"C5",x"24",x"11",x"4F",x"5F", -- 0x1F70
    x"20",x"0D",x"DC",x"CD",x"D3",x"C5",x"25",x"05", -- 0x1F78
    x"10",x"93",x"D5",x"25",x"02",x"DC",x"D5",x"DD", -- 0x1F80
    x"C5",x"0D",x"D8",x"26",x"02",x"8D",x"50",x"35", -- 0x1F88
    x"06",x"04",x"D8",x"25",x"05",x"10",x"93",x"D9", -- 0x1F90
    x"27",x"0C",x"5C",x"C1",x"08",x"26",x"04",x"4C", -- 0x1F98
    x"5F",x"84",x"07",x"7E",x"9E",x"FD",x"39",x"9E", -- 0x1FA0
    x"CF",x"EC",x"C4",x"27",x"07",x"83",x"00",x"01", -- 0x1FA8
    x"8D",x"03",x"1F",x"21",x"39",x"34",x"76",x"6F", -- 0x1FB0
    x"64",x"A6",x"63",x"3D",x"ED",x"66",x"EC",x"61", -- 0x1FB8
    x"3D",x"EB",x"66",x"89",x"00",x"ED",x"65",x"E6", -- 0x1FC0
    x"E4",x"A6",x"63",x"3D",x"E3",x"65",x"ED",x"65", -- 0x1FC8
    x"24",x"02",x"6C",x"64",x"A6",x"E4",x"E6",x"62", -- 0x1FD0
    x"3D",x"E3",x"64",x"ED",x"64",x"35",x"F6",x"7E", -- 0x1FD8
    x"94",x"A1",x"5F",x"9D",x"A5",x"27",x"11",x"BD", -- 0x1FE0
    x"B2",x"6D",x"BD",x"B1",x"41",x"96",x"4F",x"8B", -- 0x1FE8
    x"06",x"97",x"4F",x"BD",x"B7",x"0E",x"C4",x"3F", -- 0x1FF0
    x"1F",x"98",x"C4",x"07",x"44",x"44",x"44",x"39", -- 0x1FF8
    x"A1",x"CB",x"A2",x"82",x"A7",x"7C",x"A7",x"0B", -- 0x2000
    x"A7",x"F4",x"A9",x"DE",x"A7",x"D8",x"10",x"CE", -- 0x2008
    x"03",x"D7",x"86",x"37",x"B7",x"FF",x"23",x"96", -- 0x2010
    x"71",x"81",x"55",x"26",x"57",x"9E",x"72",x"A6", -- 0x2018
    x"84",x"81",x"12",x"26",x"4F",x"6E",x"84",x"31", -- 0x2020
    x"8C",x"E4",x"86",x"3A",x"B7",x"FF",x"A2",x"8E", -- 0x2028
    x"FF",x"20",x"CC",x"FF",x"34",x"6F",x"01",x"6F", -- 0x2030
    x"03",x"4A",x"A7",x"84",x"86",x"F8",x"A7",x"02", -- 0x2038
    x"E7",x"01",x"E7",x"03",x"6F",x"02",x"86",x"02", -- 0x2040
    x"A7",x"84",x"86",x"FF",x"8E",x"FF",x"00",x"6F", -- 0x2048
    x"01",x"6F",x"03",x"6F",x"84",x"A7",x"02",x"E7", -- 0x2050
    x"01",x"E7",x"03",x"7E",x"A0",x"72",x"BD",x"8C", -- 0x2058
    x"2E",x"7E",x"C0",x"00",x"E5",x"02",x"27",x"0A", -- 0x2060
    x"6F",x"1E",x"E5",x"02",x"27",x"02",x"33",x"5E", -- 0x2068
    x"A7",x"5D",x"6E",x"A4",x"8E",x"04",x"01",x"6F", -- 0x2070
    x"83",x"30",x"01",x"26",x"FA",x"BD",x"A9",x"28", -- 0x2078
    x"6F",x"80",x"9F",x"19",x"8E",x"7F",x"FF",x"20", -- 0x2080
    x"0A",x"12",x"12",x"12",x"12",x"12",x"12",x"12", -- 0x2088
    x"12",x"12",x"12",x"9F",x"74",x"9F",x"27",x"9F", -- 0x2090
    x"23",x"30",x"89",x"FF",x"38",x"9F",x"21",x"1F", -- 0x2098
    x"14",x"8E",x"A1",x"0D",x"CE",x"00",x"8F",x"C6", -- 0x20A0
    x"1C",x"BD",x"A5",x"9A",x"CE",x"01",x"0C",x"C6", -- 0x20A8
    x"1E",x"BD",x"A5",x"9A",x"AE",x"14",x"AF",x"43", -- 0x20B0
    x"AF",x"48",x"8E",x"01",x"5E",x"CC",x"39",x"4B", -- 0x20B8
    x"A7",x"80",x"5A",x"26",x"FB",x"B7",x"02",x"D9", -- 0x20C0
    x"BD",x"AD",x"19",x"7E",x"80",x"02",x"34",x"14", -- 0x20C8
    x"0D",x"E7",x"10",x"26",x"56",x"A8",x"BD",x"A1", -- 0x20D0
    x"99",x"BD",x"A1",x"CB",x"27",x"F8",x"7E",x"A1", -- 0x20D8
    x"B9",x"72",x"86",x"55",x"97",x"71",x"20",x"0B", -- 0x20E0
    x"12",x"0F",x"6F",x"BD",x"AD",x"33",x"1C",x"AF", -- 0x20E8
    x"BD",x"A9",x"10",x"7E",x"AC",x"73",x"7D",x"FF", -- 0x20F0
    x"23",x"2B",x"01",x"3B",x"BD",x"8C",x"28",x"BD", -- 0x20F8
    x"A7",x"D1",x"31",x"8C",x"03",x"7E",x"A0",x"2A", -- 0x2100
    x"0F",x"71",x"7E",x"C0",x"00",x"12",x"18",x"0A", -- 0x2108
    x"00",x"80",x"0B",x"00",x"58",x"00",x"01",x"10", -- 0x2110
    x"70",x"84",x"00",x"B4",x"4A",x"0C",x"A7",x"26", -- 0x2118
    x"02",x"0C",x"A6",x"B6",x"00",x"00",x"7E",x"AA", -- 0x2120
    x"1A",x"7E",x"A9",x"B3",x"7E",x"A0",x"F6",x"7E", -- 0x2128
    x"B4",x"4A",x"80",x"4F",x"C7",x"52",x"59",x"FF", -- 0x2130
    x"04",x"5E",x"7E",x"B2",x"77",x"35",x"AA",x"66", -- 0x2138
    x"AB",x"67",x"14",x"AB",x"1A",x"AA",x"29",x"43", -- 0x2140
    x"4F",x"4C",x"4F",x"52",x"20",x"42",x"41",x"53", -- 0x2148
    x"49",x"43",x"20",x"31",x"2E",x"32",x"0D",x"28", -- 0x2150
    x"43",x"29",x"20",x"31",x"39",x"38",x"32",x"20", -- 0x2158
    x"54",x"41",x"4E",x"44",x"59",x"00",x"4D",x"49", -- 0x2160
    x"43",x"52",x"4F",x"53",x"4F",x"46",x"54",x"0D", -- 0x2168
    x"00",x"8D",x"03",x"84",x"7F",x"39",x"BD",x"01", -- 0x2170
    x"6A",x"0F",x"70",x"0D",x"6F",x"27",x"32",x"0D", -- 0x2178
    x"79",x"26",x"03",x"03",x"70",x"39",x"34",x"74", -- 0x2180
    x"9E",x"7A",x"A6",x"80",x"34",x"02",x"9F",x"7A", -- 0x2188
    x"0A",x"79",x"26",x"03",x"BD",x"A6",x"35",x"35", -- 0x2190
    x"F6",x"0A",x"94",x"26",x"0E",x"C6",x"0B",x"D7", -- 0x2198
    x"94",x"9E",x"88",x"A6",x"84",x"8B",x"10",x"8A", -- 0x21A0
    x"8F",x"A7",x"84",x"8E",x"04",x"5E",x"7E",x"A7", -- 0x21A8
    x"D3",x"34",x"14",x"8D",x"E4",x"8D",x"14",x"27", -- 0x21B0
    x"FA",x"C6",x"60",x"E7",x"9F",x"00",x"88",x"35", -- 0x21B8
    x"94",x"7E",x"A1",x"CB",x"39",x"39",x"39",x"39", -- 0x21C0
    x"39",x"39",x"39",x"34",x"54",x"CE",x"FF",x"00", -- 0x21C8
    x"8E",x"01",x"52",x"4F",x"4A",x"34",x"12",x"A7", -- 0x21D0
    x"42",x"69",x"42",x"24",x"43",x"6C",x"60",x"8D", -- 0x21D8
    x"59",x"A7",x"61",x"A8",x"84",x"A4",x"84",x"E6", -- 0x21E0
    x"61",x"E7",x"80",x"4D",x"27",x"EB",x"E6",x"42", -- 0x21E8
    x"E7",x"62",x"C6",x"F8",x"CB",x"08",x"44",x"24", -- 0x21F0
    x"FB",x"EB",x"60",x"27",x"48",x"C1",x"1A",x"22", -- 0x21F8
    x"46",x"CA",x"40",x"8D",x"29",x"BA",x"01",x"1A", -- 0x2200
    x"26",x"02",x"CA",x"20",x"E7",x"60",x"BE",x"01", -- 0x2208
    x"1B",x"8D",x"9B",x"C6",x"FF",x"8D",x"21",x"4C", -- 0x2210
    x"26",x"06",x"E6",x"62",x"8D",x"1A",x"A1",x"61", -- 0x2218
    x"35",x"12",x"26",x"07",x"81",x"12",x"26",x"04", -- 0x2220
    x"73",x"01",x"1A",x"4F",x"35",x"D4",x"86",x"7F", -- 0x2228
    x"A7",x"42",x"A6",x"C4",x"43",x"84",x"40",x"39", -- 0x2230
    x"E7",x"42",x"A6",x"C4",x"8A",x"80",x"6D",x"42", -- 0x2238
    x"2B",x"02",x"8A",x"C0",x"39",x"C6",x"33",x"8E", -- 0x2240
    x"A2",x"38",x"C1",x"21",x"25",x"16",x"8E",x"A2", -- 0x2248
    x"1A",x"C1",x"30",x"24",x"0F",x"8D",x"D7",x"C1", -- 0x2250
    x"2B",x"23",x"02",x"88",x"40",x"4D",x"26",x"AC", -- 0x2258
    x"CB",x"10",x"20",x"A8",x"58",x"8D",x"C7",x"27", -- 0x2260
    x"01",x"5C",x"E6",x"85",x"20",x"9E",x"5E",x"5F", -- 0x2268
    x"0A",x"5B",x"08",x"15",x"09",x"5D",x"20",x"20", -- 0x2270
    x"30",x"12",x"0D",x"0D",x"0C",x"5C",x"03",x"03", -- 0x2278
    x"40",x"13",x"BD",x"01",x"67",x"34",x"04",x"D6", -- 0x2280
    x"6F",x"5C",x"35",x"04",x"2B",x"31",x"26",x"7A", -- 0x2288
    x"34",x"16",x"D6",x"78",x"5A",x"27",x"0F",x"D6", -- 0x2290
    x"79",x"5C",x"26",x"02",x"8D",x"0A",x"9E",x"7A", -- 0x2298
    x"A7",x"80",x"9F",x"7A",x"0C",x"79",x"35",x"96", -- 0x22A0
    x"C6",x"01",x"D7",x"7C",x"8E",x"01",x"DA",x"9F", -- 0x22A8
    x"7E",x"D6",x"79",x"D7",x"7D",x"34",x"62",x"BD", -- 0x22B0
    x"A7",x"E5",x"35",x"62",x"7E",x"A6",x"50",x"34", -- 0x22B8
    x"17",x"1A",x"50",x"F6",x"FF",x"22",x"54",x"25", -- 0x22C0
    x"FA",x"8D",x"30",x"5F",x"8D",x"2F",x"C6",x"08", -- 0x22C8
    x"34",x"04",x"5F",x"44",x"59",x"58",x"8D",x"25", -- 0x22D0
    x"35",x"04",x"5A",x"26",x"F3",x"8D",x"1C",x"35", -- 0x22D8
    x"03",x"81",x"0D",x"27",x"08",x"0C",x"9C",x"D6", -- 0x22E0
    x"9C",x"D1",x"9B",x"25",x"06",x"0F",x"9C",x"8D", -- 0x22E8
    x"14",x"8D",x"12",x"F6",x"FF",x"22",x"54",x"25", -- 0x22F0
    x"FA",x"35",x"94",x"C6",x"02",x"F7",x"FF",x"20", -- 0x22F8
    x"8D",x"00",x"9E",x"95",x"8C",x"9E",x"97",x"7E", -- 0x2300
    x"A7",x"D3",x"34",x"16",x"9E",x"88",x"81",x"08", -- 0x2308
    x"26",x"0B",x"8C",x"04",x"00",x"27",x"46",x"86", -- 0x2310
    x"60",x"A7",x"82",x"20",x"27",x"81",x"0D",x"26", -- 0x2318
    x"0E",x"9E",x"88",x"86",x"60",x"A7",x"80",x"1F", -- 0x2320
    x"10",x"C5",x"1F",x"26",x"F6",x"20",x"15",x"81", -- 0x2328
    x"20",x"25",x"2A",x"4D",x"2B",x"0C",x"81",x"40", -- 0x2330
    x"25",x"06",x"81",x"60",x"25",x"04",x"84",x"DF", -- 0x2338
    x"88",x"40",x"A7",x"80",x"9F",x"88",x"8C",x"05", -- 0x2340
    x"FF",x"23",x"12",x"8E",x"04",x"00",x"EC",x"88", -- 0x2348
    x"20",x"ED",x"81",x"8C",x"05",x"E0",x"25",x"F6", -- 0x2350
    x"C6",x"60",x"BD",x"A9",x"2D",x"35",x"96",x"BD", -- 0x2358
    x"01",x"64",x"34",x"16",x"0F",x"6E",x"96",x"6F", -- 0x2360
    x"27",x"09",x"4C",x"27",x"17",x"9E",x"99",x"DC", -- 0x2368
    x"9B",x"20",x"09",x"D6",x"89",x"C4",x"1F",x"8E", -- 0x2370
    x"10",x"10",x"86",x"20",x"9F",x"6A",x"D7",x"6C", -- 0x2378
    x"97",x"6D",x"35",x"96",x"03",x"6E",x"8E",x"01", -- 0x2380
    x"00",x"4F",x"5F",x"20",x"EF",x"BD",x"A9",x"28", -- 0x2388
    x"BD",x"01",x"82",x"0F",x"87",x"8E",x"02",x"DD", -- 0x2390
    x"C6",x"01",x"BD",x"A1",x"71",x"0D",x"70",x"26", -- 0x2398
    x"2B",x"0D",x"6F",x"26",x"23",x"81",x"0C",x"27", -- 0x23A0
    x"E4",x"81",x"08",x"26",x"07",x"5A",x"27",x"E0", -- 0x23A8
    x"30",x"1F",x"20",x"34",x"81",x"15",x"26",x"0A", -- 0x23B0
    x"5A",x"27",x"D5",x"86",x"08",x"BD",x"A2",x"82", -- 0x23B8
    x"20",x"F6",x"81",x"03",x"1A",x"01",x"27",x"05", -- 0x23C0
    x"81",x"0D",x"26",x"0D",x"4F",x"34",x"01",x"BD", -- 0x23C8
    x"B9",x"58",x"6F",x"84",x"8E",x"02",x"DC",x"35", -- 0x23D0
    x"81",x"81",x"20",x"25",x"BD",x"81",x"7B",x"24", -- 0x23D8
    x"B9",x"C1",x"FA",x"24",x"B5",x"A7",x"80",x"5C", -- 0x23E0
    x"BD",x"A2",x"82",x"20",x"AD",x"BD",x"01",x"6D", -- 0x23E8
    x"96",x"6F",x"27",x"21",x"4C",x"26",x"0C",x"96", -- 0x23F0
    x"78",x"26",x"05",x"C6",x"2C",x"7E",x"AC",x"46", -- 0x23F8
    x"4A",x"27",x"12",x"7E",x"A6",x"16",x"BD",x"01", -- 0x2400
    x"70",x"96",x"6F",x"4C",x"26",x"07",x"96",x"78", -- 0x2408
    x"27",x"E9",x"4A",x"27",x"EE",x"39",x"27",x"0E", -- 0x2410
    x"BD",x"A5",x"A5",x"8D",x"10",x"9D",x"A5",x"27", -- 0x2418
    x"2A",x"BD",x"A5",x"A2",x"20",x"F5",x"BD",x"01", -- 0x2420
    x"73",x"86",x"FF",x"97",x"6F",x"BD",x"01",x"76", -- 0x2428
    x"96",x"6F",x"0F",x"6F",x"4C",x"26",x"14",x"96", -- 0x2430
    x"78",x"81",x"02",x"26",x"0C",x"96",x"79",x"27", -- 0x2438
    x"03",x"BD",x"A2",x"A8",x"C6",x"FF",x"BD",x"A2", -- 0x2440
    x"AA",x"0F",x"78",x"39",x"BD",x"A5",x"78",x"9D", -- 0x2448
    x"A5",x"27",x"16",x"BD",x"B2",x"6D",x"C6",x"41", -- 0x2450
    x"BD",x"B2",x"6F",x"26",x"EE",x"4F",x"BD",x"A6", -- 0x2458
    x"5C",x"86",x"FF",x"97",x"6F",x"4F",x"7E",x"B7", -- 0x2460
    x"64",x"4F",x"9E",x"8A",x"BD",x"A6",x"5F",x"0F", -- 0x2468
    x"78",x"0C",x"7C",x"BD",x"A7",x"D8",x"9E",x"19", -- 0x2470
    x"9F",x"7E",x"86",x"FF",x"97",x"7D",x"DC",x"1B", -- 0x2478
    x"93",x"7E",x"27",x"0D",x"10",x"83",x"00",x"FF", -- 0x2480
    x"24",x"02",x"D7",x"7D",x"BD",x"A7",x"F4",x"20", -- 0x2488
    x"E7",x"00",x"7C",x"0F",x"7D",x"7E",x"A7",x"E7", -- 0x2490
    x"0F",x"78",x"81",x"4D",x"27",x"60",x"32",x"62", -- 0x2498
    x"BD",x"A5",x"C5",x"BD",x"A6",x"48",x"7D",x"01", -- 0x24A0
    x"E4",x"27",x"1D",x"B6",x"01",x"E3",x"27",x"1D", -- 0x24A8
    x"BD",x"AD",x"19",x"86",x"FF",x"97",x"6F",x"0C", -- 0x24B0
    x"78",x"BD",x"A6",x"35",x"7E",x"AC",x"7C",x"BD", -- 0x24B8
    x"01",x"85",x"BD",x"A4",x"2D",x"7E",x"AC",x"73", -- 0x24C0
    x"B6",x"01",x"E2",x"27",x"03",x"7E",x"A6",x"16", -- 0x24C8
    x"BD",x"AD",x"19",x"BD",x"A7",x"7C",x"9E",x"19", -- 0x24D0
    x"9F",x"7E",x"DC",x"7E",x"4C",x"BD",x"AC",x"37", -- 0x24D8
    x"BD",x"A7",x"0B",x"26",x"13",x"96",x"7C",x"27", -- 0x24E0
    x"0F",x"2A",x"ED",x"9F",x"1B",x"8D",x"4C",x"8E", -- 0x24E8
    x"AB",x"EC",x"BD",x"B9",x"9C",x"7E",x"AC",x"E9", -- 0x24F0
    x"BD",x"AD",x"19",x"7E",x"A6",x"19",x"9D",x"9F", -- 0x24F8
    x"8D",x"76",x"BD",x"A6",x"48",x"9E",x"8A",x"9D", -- 0x2500
    x"A5",x"27",x"06",x"BD",x"B2",x"6D",x"BD",x"B7", -- 0x2508
    x"3D",x"B6",x"01",x"E2",x"81",x"02",x"26",x"B5", -- 0x2510
    x"FC",x"01",x"E5",x"33",x"8B",x"DF",x"9D",x"7D", -- 0x2518
    x"01",x"E4",x"26",x"A9",x"FC",x"01",x"E7",x"30", -- 0x2520
    x"8B",x"9F",x"7E",x"BD",x"A7",x"7C",x"BD",x"A7", -- 0x2528
    x"0B",x"26",x"C8",x"9F",x"7E",x"0D",x"7C",x"27", -- 0x2530
    x"C2",x"2A",x"F3",x"7E",x"A7",x"E9",x"27",x"05", -- 0x2538
    x"BD",x"B7",x"3D",x"9F",x"9D",x"6E",x"9F",x"00", -- 0x2540
    x"9D",x"BD",x"01",x"7F",x"96",x"6F",x"4C",x"27", -- 0x2548
    x"50",x"7E",x"AD",x"EB",x"BD",x"B3",x"E4",x"83", -- 0x2550
    x"01",x"FF",x"10",x"22",x"0E",x"EC",x"C3",x"05", -- 0x2558
    x"FF",x"DD",x"88",x"39",x"96",x"87",x"26",x"03", -- 0x2560
    x"BD",x"A1",x"CB",x"0F",x"87",x"97",x"53",x"10", -- 0x2568
    x"26",x"11",x"1C",x"97",x"56",x"7E",x"B6",x"9B", -- 0x2570
    x"8E",x"01",x"D1",x"6F",x"80",x"86",x"20",x"A7", -- 0x2578
    x"80",x"8C",x"01",x"DA",x"26",x"F9",x"9D",x"A5", -- 0x2580
    x"27",x"17",x"BD",x"B1",x"56",x"BD",x"B6",x"54", -- 0x2588
    x"CE",x"01",x"D1",x"E7",x"C0",x"27",x"0A",x"8C", -- 0x2590
    x"C6",x"08",x"A6",x"80",x"A7",x"C0",x"5A",x"26", -- 0x2598
    x"F9",x"39",x"BD",x"B2",x"6D",x"81",x"23",x"26", -- 0x25A0
    x"02",x"9D",x"9F",x"BD",x"B1",x"41",x"BD",x"B3", -- 0x25A8
    x"ED",x"59",x"89",x"00",x"26",x"69",x"56",x"D7", -- 0x25B0
    x"6F",x"BD",x"01",x"61",x"27",x"06",x"2A",x"5F", -- 0x25B8
    x"C1",x"FE",x"2D",x"5B",x"39",x"8D",x"B1",x"9D", -- 0x25C0
    x"A5",x"27",x"F9",x"7E",x"B2",x"77",x"BD",x"01", -- 0x25C8
    x"88",x"96",x"6F",x"34",x"02",x"8D",x"D7",x"BD", -- 0x25D0
    x"A3",x"ED",x"5F",x"96",x"6F",x"27",x"05",x"0D", -- 0x25D8
    x"79",x"26",x"01",x"53",x"35",x"02",x"97",x"6F", -- 0x25E0
    x"1D",x"7E",x"B4",x"F4",x"8D",x"D7",x"8D",x"58", -- 0x25E8
    x"BD",x"A6",x"D1",x"26",x"24",x"39",x"BD",x"01", -- 0x25F0
    x"5E",x"BD",x"B1",x"56",x"BD",x"B6",x"A4",x"34", -- 0x25F8
    x"04",x"8D",x"9F",x"BD",x"B2",x"6D",x"8D",x"BD", -- 0x2600
    x"96",x"6F",x"0F",x"6F",x"35",x"04",x"C1",x"49", -- 0x2608
    x"27",x"12",x"C1",x"4F",x"27",x"42",x"C6",x"2A", -- 0x2610
    x"8C",x"C6",x"28",x"8C",x"C6",x"24",x"8C",x"C6", -- 0x2618
    x"26",x"7E",x"AC",x"46",x"4C",x"2B",x"EF",x"26", -- 0x2620
    x"2E",x"8D",x"1D",x"B6",x"01",x"E3",x"B4",x"01", -- 0x2628
    x"E4",x"27",x"E3",x"0C",x"78",x"BD",x"A7",x"01", -- 0x2630
    x"26",x"DF",x"0D",x"7C",x"27",x"DB",x"2B",x"17", -- 0x2638
    x"96",x"7D",x"27",x"F1",x"97",x"79",x"20",x"0A", -- 0x2640
    x"0D",x"78",x"26",x"D0",x"8D",x"33",x"26",x"C9", -- 0x2648
    x"0F",x"79",x"8E",x"01",x"DA",x"9F",x"7A",x"39", -- 0x2650
    x"4C",x"26",x"FC",x"4C",x"8E",x"FF",x"FF",x"0D", -- 0x2658
    x"78",x"26",x"B9",x"CE",x"01",x"DA",x"DF",x"7E", -- 0x2660
    x"A7",x"48",x"AF",x"49",x"8E",x"01",x"D2",x"BD", -- 0x2668
    x"A5",x"98",x"0F",x"7C",x"86",x"0F",x"97",x"7D", -- 0x2670
    x"BD",x"A7",x"E5",x"86",x"02",x"97",x"78",x"20", -- 0x2678
    x"CF",x"8E",x"01",x"DA",x"9F",x"7E",x"96",x"68", -- 0x2680
    x"4C",x"26",x"0B",x"BD",x"A9",x"28",x"9E",x"88", -- 0x2688
    x"C6",x"53",x"E7",x"81",x"9F",x"88",x"8D",x"69", -- 0x2690
    x"DA",x"7C",x"26",x"34",x"8E",x"01",x"DA",x"CE", -- 0x2698
    x"01",x"D2",x"C6",x"08",x"6F",x"E2",x"A6",x"80", -- 0x26A0
    x"10",x"9E",x"68",x"31",x"21",x"26",x"05",x"0F", -- 0x26A8
    x"6F",x"BD",x"A2",x"82",x"A0",x"C0",x"AA",x"E4", -- 0x26B0
    x"A7",x"E4",x"5A",x"26",x"E9",x"A6",x"E0",x"27", -- 0x26B8
    x"0A",x"6D",x"57",x"27",x"06",x"8D",x"0A",x"26", -- 0x26C0
    x"07",x"20",x"BB",x"86",x"46",x"8D",x"29",x"4F", -- 0x26C8
    x"39",x"7D",x"01",x"E4",x"26",x"09",x"BD",x"A7", -- 0x26D0
    x"7C",x"8D",x"30",x"8D",x"08",x"20",x"FA",x"8D", -- 0x26D8
    x"20",x"8D",x"02",x"20",x"FA",x"26",x"06",x"96", -- 0x26E0
    x"7C",x"40",x"2B",x"14",x"4A",x"97",x"81",x"32", -- 0x26E8
    x"62",x"20",x"12",x"B6",x"04",x"00",x"88",x"40", -- 0x26F0
    x"D6",x"68",x"5C",x"26",x"03",x"B7",x"04",x"00", -- 0x26F8
    x"39",x"8D",x"79",x"8D",x"06",x"BD",x"A7",x"E9", -- 0x2700
    x"D6",x"81",x"39",x"1A",x"50",x"8D",x"E4",x"9E", -- 0x2708
    x"7E",x"4F",x"8D",x"41",x"46",x"81",x"3C",x"26", -- 0x2710
    x"F9",x"8D",x"2E",x"97",x"7C",x"8D",x"2A",x"97", -- 0x2718
    x"7D",x"9B",x"7C",x"97",x"80",x"96",x"7D",x"97", -- 0x2720
    x"81",x"27",x"10",x"8D",x"1C",x"A7",x"84",x"A1", -- 0x2728
    x"80",x"26",x"11",x"9B",x"80",x"97",x"80",x"0A", -- 0x2730
    x"81",x"26",x"F0",x"8D",x"0C",x"90",x"80",x"27", -- 0x2738
    x"05",x"86",x"01",x"8C",x"86",x"02",x"97",x"81", -- 0x2740
    x"39",x"86",x"08",x"97",x"82",x"8D",x"06",x"46", -- 0x2748
    x"0A",x"82",x"26",x"F9",x"39",x"8D",x"06",x"D6", -- 0x2750
    x"83",x"5A",x"D1",x"8F",x"39",x"0F",x"83",x"0D", -- 0x2758
    x"84",x"26",x"10",x"8D",x"07",x"25",x"FC",x"8D", -- 0x2760
    x"03",x"24",x"FC",x"39",x"0C",x"83",x"F6",x"FF", -- 0x2768
    x"20",x"56",x"39",x"8D",x"F7",x"24",x"FC",x"8D", -- 0x2770
    x"F3",x"25",x"FC",x"39",x"1A",x"50",x"8D",x"4A", -- 0x2778
    x"0F",x"82",x"8D",x"DF",x"8D",x"27",x"22",x"0F", -- 0x2780
    x"8D",x"1D",x"25",x"0F",x"0A",x"82",x"96",x"82", -- 0x2788
    x"81",x"A0",x"26",x"EE",x"97",x"84",x"39",x"8D", -- 0x2790
    x"0E",x"22",x"E9",x"8D",x"10",x"25",x"E9",x"0C", -- 0x2798
    x"82",x"96",x"82",x"80",x"60",x"20",x"EB",x"0F", -- 0x27A0
    x"83",x"8D",x"BC",x"20",x"04",x"0F",x"83",x"8D", -- 0x27A8
    x"C6",x"D6",x"83",x"D1",x"90",x"22",x"03",x"D1", -- 0x27B0
    x"91",x"39",x"0F",x"82",x"39",x"1F",x"89",x"9D", -- 0x27B8
    x"9F",x"C1",x"AA",x"27",x"24",x"C1",x"88",x"BD", -- 0x27C0
    x"A5",x"C9",x"B6",x"FF",x"21",x"8A",x"08",x"8D", -- 0x27C8
    x"1F",x"9E",x"8A",x"30",x"1F",x"26",x"FC",x"39", -- 0x27D0
    x"1A",x"50",x"8D",x"EE",x"9E",x"92",x"8D",x"48", -- 0x27D8
    x"30",x"1F",x"26",x"FA",x"39",x"8D",x"F1",x"8D", -- 0x27E0
    x"0B",x"1C",x"AF",x"B6",x"FF",x"21",x"84",x"F7", -- 0x27E8
    x"B7",x"FF",x"21",x"39",x"1A",x"50",x"D6",x"7D", -- 0x27F0
    x"D7",x"81",x"96",x"7D",x"27",x"07",x"9E",x"7E", -- 0x27F8
    x"AB",x"80",x"5A",x"26",x"FB",x"9B",x"7C",x"97", -- 0x2800
    x"80",x"9E",x"7E",x"8D",x"1B",x"86",x"3C",x"8D", -- 0x2808
    x"19",x"96",x"7C",x"8D",x"15",x"96",x"7D",x"8D", -- 0x2810
    x"11",x"4D",x"27",x"08",x"A6",x"80",x"8D",x"0A", -- 0x2818
    x"0A",x"81",x"26",x"F8",x"96",x"80",x"8D",x"02", -- 0x2820
    x"86",x"55",x"34",x"02",x"C6",x"01",x"96",x"85", -- 0x2828
    x"B7",x"FF",x"20",x"10",x"8E",x"A8",x"5C",x"E5", -- 0x2830
    x"E4",x"26",x"0D",x"A6",x"A0",x"10",x"8C",x"A8", -- 0x2838
    x"80",x"27",x"12",x"B7",x"FF",x"20",x"20",x"F3", -- 0x2840
    x"A6",x"A1",x"10",x"8C",x"A8",x"80",x"27",x"05", -- 0x2848
    x"B7",x"FF",x"20",x"20",x"F3",x"97",x"85",x"58", -- 0x2850
    x"24",x"D4",x"35",x"82",x"82",x"92",x"AA",x"BA", -- 0x2858
    x"CA",x"DA",x"EA",x"F2",x"FA",x"FA",x"FA",x"F2", -- 0x2860
    x"EA",x"DA",x"CA",x"BA",x"AA",x"92",x"7A",x"6A", -- 0x2868
    x"52",x"42",x"32",x"22",x"12",x"0A",x"02",x"02", -- 0x2870
    x"02",x"0A",x"12",x"22",x"32",x"42",x"52",x"6A", -- 0x2878
    x"8D",x"3F",x"34",x"10",x"BD",x"B7",x"38",x"35", -- 0x2880
    x"10",x"C1",x"08",x"22",x"48",x"5A",x"2B",x"05", -- 0x2888
    x"86",x"10",x"3D",x"20",x"08",x"E6",x"84",x"2A", -- 0x2890
    x"03",x"C4",x"70",x"21",x"5F",x"34",x"04",x"8D", -- 0x2898
    x"6C",x"A6",x"84",x"2B",x"01",x"4F",x"84",x"0F", -- 0x28A0
    x"9A",x"86",x"AA",x"E0",x"8A",x"80",x"A7",x"84", -- 0x28A8
    x"39",x"8D",x"0E",x"8D",x"58",x"4F",x"E6",x"84", -- 0x28B0
    x"2A",x"F2",x"03",x"86",x"D4",x"86",x"E7",x"84", -- 0x28B8
    x"39",x"BD",x"B2",x"6A",x"BD",x"01",x"9D",x"BD", -- 0x28C0
    x"B7",x"0B",x"C1",x"3F",x"22",x"07",x"34",x"04", -- 0x28C8
    x"BD",x"B7",x"38",x"C1",x"1F",x"22",x"71",x"34", -- 0x28D0
    x"04",x"54",x"86",x"20",x"3D",x"8E",x"04",x"00", -- 0x28D8
    x"30",x"8B",x"E6",x"61",x"54",x"3A",x"35",x"06", -- 0x28E0
    x"84",x"01",x"56",x"49",x"C6",x"10",x"54",x"4A", -- 0x28E8
    x"2A",x"FC",x"D7",x"86",x"39",x"8D",x"CD",x"C6", -- 0x28F0
    x"FF",x"A6",x"84",x"2A",x"0D",x"94",x"86",x"27", -- 0x28F8
    x"08",x"E6",x"84",x"54",x"54",x"54",x"54",x"C4", -- 0x2900
    x"07",x"5C",x"BD",x"A5",x"E8",x"7E",x"B2",x"67", -- 0x2908
    x"BD",x"01",x"A0",x"27",x"13",x"BD",x"B7",x"0B", -- 0x2910
    x"C1",x"08",x"22",x"1B",x"5D",x"27",x"06",x"5A", -- 0x2918
    x"86",x"10",x"3D",x"CA",x"0F",x"CA",x"80",x"8C", -- 0x2920
    x"C6",x"60",x"8E",x"04",x"00",x"9F",x"88",x"E7", -- 0x2928
    x"80",x"8C",x"05",x"FF",x"23",x"F9",x"39",x"8D", -- 0x2930
    x"EF",x"8E",x"A1",x"65",x"7E",x"B9",x"9C",x"BD", -- 0x2938
    x"B2",x"6D",x"BD",x"B7",x"0B",x"5D",x"26",x"3C", -- 0x2940
    x"7E",x"B4",x"4A",x"8D",x"F5",x"D7",x"8C",x"8D", -- 0x2948
    x"EE",x"86",x"04",x"3D",x"DD",x"8D",x"B6",x"FF", -- 0x2950
    x"03",x"8A",x"01",x"B7",x"FF",x"03",x"0F",x"08", -- 0x2958
    x"8D",x"40",x"8D",x"12",x"8D",x"1F",x"86",x"FE", -- 0x2960
    x"8D",x"1D",x"8D",x"19",x"86",x"02",x"8D",x"17", -- 0x2968
    x"9E",x"8D",x"26",x"F0",x"4F",x"8C",x"86",x"08", -- 0x2970
    x"A7",x"E2",x"B6",x"FF",x"23",x"84",x"F7",x"AA", -- 0x2978
    x"E0",x"B7",x"FF",x"23",x"39",x"86",x"7E",x"B7", -- 0x2980
    x"FF",x"20",x"96",x"8C",x"4C",x"26",x"FD",x"39", -- 0x2988
    x"1F",x"89",x"9D",x"9F",x"C1",x"AA",x"27",x"DC", -- 0x2990
    x"C0",x"88",x"BD",x"A5",x"C9",x"5C",x"8D",x"02", -- 0x2998
    x"20",x"D4",x"CE",x"FF",x"01",x"8D",x"00",x"A6", -- 0x29A0
    x"C4",x"84",x"F7",x"57",x"24",x"02",x"8A",x"08", -- 0x29A8
    x"A7",x"C1",x"39",x"B6",x"FF",x"03",x"2A",x"0D", -- 0x29B0
    x"B6",x"FF",x"02",x"BE",x"00",x"8D",x"27",x"05", -- 0x29B8
    x"30",x"1F",x"BF",x"00",x"8D",x"3B",x"BD",x"B7", -- 0x29C0
    x"0E",x"C1",x"03",x"10",x"22",x"0A",x"7B",x"5D", -- 0x29C8
    x"26",x"02",x"8D",x"0A",x"8E",x"01",x"5A",x"D6", -- 0x29D0
    x"53",x"E6",x"85",x"7E",x"B4",x"F3",x"8D",x"94", -- 0x29D8
    x"8E",x"01",x"5E",x"C6",x"03",x"86",x"0A",x"ED", -- 0x29E0
    x"E3",x"8D",x"B7",x"CC",x"40",x"80",x"A7",x"E2", -- 0x29E8
    x"CA",x"02",x"F7",x"FF",x"20",x"C8",x"02",x"B6", -- 0x29F0
    x"FF",x"00",x"2B",x"03",x"E0",x"E4",x"8C",x"EB", -- 0x29F8
    x"E4",x"A6",x"E0",x"44",x"81",x"01",x"26",x"E6", -- 0x2A00
    x"54",x"54",x"E1",x"1F",x"27",x"04",x"6A",x"E4", -- 0x2A08
    x"26",x"D9",x"E7",x"82",x"EC",x"E1",x"5A",x"2A", -- 0x2A10
    x"CC",x"39",x"81",x"3A",x"24",x"0A",x"81",x"20", -- 0x2A18
    x"26",x"02",x"0E",x"9F",x"80",x"30",x"80",x"D0", -- 0x2A20
    x"39",x"BC",x"7A",x"BC",x"EE",x"BC",x"93",x"01", -- 0x2A28
    x"12",x"BF",x"1F",x"BF",x"78",x"B7",x"50",x"B6", -- 0x2A30
    x"81",x"B4",x"FD",x"B7",x"16",x"B6",x"A0",x"B6", -- 0x2A38
    x"8C",x"A5",x"CE",x"A9",x"C6",x"B6",x"AB",x"B6", -- 0x2A40
    x"C8",x"B6",x"CF",x"A8",x"F5",x"A5",x"64",x"B4", -- 0x2A48
    x"EE",x"79",x"B9",x"C5",x"79",x"B9",x"BC",x"7B", -- 0x2A50
    x"BA",x"CC",x"7B",x"BB",x"91",x"7F",x"01",x"1D", -- 0x2A58
    x"50",x"B2",x"D5",x"46",x"B2",x"D4",x"46",x"4F", -- 0x2A60
    x"D2",x"47",x"CF",x"52",x"45",x"CD",x"A7",x"45", -- 0x2A68
    x"4C",x"53",x"C5",x"49",x"C6",x"44",x"41",x"54", -- 0x2A70
    x"C1",x"50",x"52",x"49",x"4E",x"D4",x"4F",x"CE", -- 0x2A78
    x"49",x"4E",x"50",x"55",x"D4",x"45",x"4E",x"C4", -- 0x2A80
    x"4E",x"45",x"58",x"D4",x"44",x"49",x"CD",x"52", -- 0x2A88
    x"45",x"41",x"C4",x"52",x"55",x"CE",x"52",x"45", -- 0x2A90
    x"53",x"54",x"4F",x"52",x"C5",x"52",x"45",x"54", -- 0x2A98
    x"55",x"52",x"CE",x"53",x"54",x"4F",x"D0",x"50", -- 0x2AA0
    x"4F",x"4B",x"C5",x"43",x"4F",x"4E",x"D4",x"4C", -- 0x2AA8
    x"49",x"53",x"D4",x"43",x"4C",x"45",x"41",x"D2", -- 0x2AB0
    x"4E",x"45",x"D7",x"43",x"4C",x"4F",x"41",x"C4", -- 0x2AB8
    x"43",x"53",x"41",x"56",x"C5",x"4F",x"50",x"45", -- 0x2AC0
    x"CE",x"43",x"4C",x"4F",x"53",x"C5",x"4C",x"4C", -- 0x2AC8
    x"49",x"53",x"D4",x"53",x"45",x"D4",x"52",x"45", -- 0x2AD0
    x"53",x"45",x"D4",x"43",x"4C",x"D3",x"4D",x"4F", -- 0x2AD8
    x"54",x"4F",x"D2",x"53",x"4F",x"55",x"4E",x"C4", -- 0x2AE0
    x"41",x"55",x"44",x"49",x"CF",x"45",x"58",x"45", -- 0x2AE8
    x"C3",x"53",x"4B",x"49",x"50",x"C6",x"54",x"41", -- 0x2AF0
    x"42",x"A8",x"54",x"CF",x"53",x"55",x"C2",x"54", -- 0x2AF8
    x"48",x"45",x"CE",x"4E",x"4F",x"D4",x"53",x"54", -- 0x2B00
    x"45",x"D0",x"4F",x"46",x"C6",x"AB",x"AD",x"AA", -- 0x2B08
    x"AF",x"DE",x"41",x"4E",x"C4",x"4F",x"D2",x"BE", -- 0x2B10
    x"BD",x"BC",x"53",x"47",x"CE",x"49",x"4E",x"D4", -- 0x2B18
    x"41",x"42",x"D3",x"55",x"53",x"D2",x"52",x"4E", -- 0x2B20
    x"C4",x"53",x"49",x"CE",x"50",x"45",x"45",x"CB", -- 0x2B28
    x"4C",x"45",x"CE",x"53",x"54",x"52",x"A4",x"56", -- 0x2B30
    x"41",x"CC",x"41",x"53",x"C3",x"43",x"48",x"52", -- 0x2B38
    x"A4",x"45",x"4F",x"C6",x"4A",x"4F",x"59",x"53", -- 0x2B40
    x"54",x"CB",x"4C",x"45",x"46",x"54",x"A4",x"52", -- 0x2B48
    x"49",x"47",x"48",x"54",x"A4",x"4D",x"49",x"44", -- 0x2B50
    x"A4",x"50",x"4F",x"49",x"4E",x"D4",x"49",x"4E", -- 0x2B58
    x"4B",x"45",x"59",x"A4",x"4D",x"45",x"CD",x"AD", -- 0x2B60
    x"47",x"AE",x"86",x"AE",x"E3",x"AE",x"E3",x"AE", -- 0x2B68
    x"E3",x"AF",x"14",x"AE",x"E0",x"B8",x"F7",x"AF", -- 0x2B70
    x"42",x"AF",x"F5",x"AE",x"02",x"B0",x"F8",x"B3", -- 0x2B78
    x"4E",x"B0",x"46",x"AE",x"75",x"AD",x"E4",x"AE", -- 0x2B80
    x"C0",x"AE",x"09",x"B7",x"57",x"AE",x"30",x"B7", -- 0x2B88
    x"64",x"AE",x"41",x"AD",x"17",x"A4",x"98",x"A4", -- 0x2B90
    x"4C",x"A5",x"F6",x"A4",x"16",x"B7",x"5E",x"A8", -- 0x2B98
    x"80",x"A8",x"B1",x"A9",x"10",x"A7",x"BD",x"A9", -- 0x2BA0
    x"4B",x"A9",x"90",x"A5",x"3E",x"A5",x"EC",x"4E", -- 0x2BA8
    x"46",x"53",x"4E",x"52",x"47",x"4F",x"44",x"46", -- 0x2BB0
    x"43",x"4F",x"56",x"4F",x"4D",x"55",x"4C",x"42", -- 0x2BB8
    x"53",x"44",x"44",x"2F",x"30",x"49",x"44",x"54", -- 0x2BC0
    x"4D",x"4F",x"53",x"4C",x"53",x"53",x"54",x"43", -- 0x2BC8
    x"4E",x"46",x"44",x"41",x"4F",x"44",x"4E",x"49", -- 0x2BD0
    x"4F",x"46",x"4D",x"4E",x"4F",x"49",x"45",x"44", -- 0x2BD8
    x"53",x"20",x"45",x"52",x"52",x"4F",x"52",x"00", -- 0x2BE0
    x"20",x"49",x"4E",x"20",x"00",x"0D",x"4F",x"4B", -- 0x2BE8
    x"0D",x"00",x"0D",x"42",x"52",x"45",x"41",x"4B", -- 0x2BF0
    x"00",x"30",x"64",x"C6",x"12",x"9F",x"0F",x"A6", -- 0x2BF8
    x"84",x"80",x"80",x"26",x"15",x"AE",x"01",x"9F", -- 0x2C00
    x"11",x"9E",x"3B",x"27",x"09",x"9C",x"11",x"27", -- 0x2C08
    x"09",x"9E",x"0F",x"3A",x"20",x"E5",x"9E",x"11", -- 0x2C10
    x"9F",x"3B",x"9E",x"0F",x"4D",x"39",x"8D",x"17", -- 0x2C18
    x"DE",x"41",x"33",x"41",x"9E",x"43",x"30",x"01", -- 0x2C20
    x"A6",x"82",x"36",x"02",x"9C",x"47",x"26",x"F8", -- 0x2C28
    x"DF",x"45",x"39",x"4F",x"58",x"D3",x"1F",x"C3", -- 0x2C30
    x"00",x"3A",x"25",x"08",x"10",x"DF",x"17",x"10", -- 0x2C38
    x"93",x"17",x"25",x"EE",x"C6",x"0C",x"BD",x"01", -- 0x2C40
    x"8E",x"BD",x"01",x"91",x"BD",x"A7",x"E9",x"BD", -- 0x2C48
    x"A9",x"74",x"BD",x"AD",x"33",x"0F",x"6F",x"BD", -- 0x2C50
    x"B9",x"5C",x"BD",x"B9",x"AF",x"8E",x"AB",x"AF", -- 0x2C58
    x"3A",x"8D",x"3D",x"8D",x"3B",x"8E",x"AB",x"E0", -- 0x2C60
    x"BD",x"B9",x"9C",x"96",x"68",x"4C",x"27",x"03", -- 0x2C68
    x"BD",x"BD",x"C5",x"BD",x"B9",x"5C",x"8E",x"AB", -- 0x2C70
    x"ED",x"BD",x"B9",x"9C",x"BD",x"A3",x"90",x"CE", -- 0x2C78
    x"FF",x"FF",x"DF",x"68",x"25",x"F6",x"0D",x"70", -- 0x2C80
    x"10",x"26",x"F8",x"33",x"9F",x"A6",x"9D",x"9F", -- 0x2C88
    x"27",x"EA",x"25",x"11",x"C6",x"30",x"0D",x"6F", -- 0x2C90
    x"26",x"AC",x"BD",x"B8",x"21",x"7E",x"AD",x"C0", -- 0x2C98
    x"A6",x"80",x"7E",x"B9",x"B1",x"BD",x"AF",x"67", -- 0x2CA0
    x"9E",x"2B",x"BF",x"02",x"DA",x"BD",x"B8",x"21", -- 0x2CA8
    x"D7",x"03",x"8D",x"4D",x"25",x"12",x"DC",x"47", -- 0x2CB0
    x"A3",x"84",x"D3",x"1B",x"DD",x"1B",x"EE",x"84", -- 0x2CB8
    x"37",x"02",x"A7",x"80",x"9C",x"1B",x"26",x"F8", -- 0x2CC0
    x"B6",x"02",x"DC",x"27",x"1C",x"DC",x"1B",x"DD", -- 0x2CC8
    x"43",x"DB",x"03",x"89",x"00",x"DD",x"41",x"BD", -- 0x2CD0
    x"AC",x"1E",x"CE",x"02",x"D8",x"37",x"02",x"A7", -- 0x2CD8
    x"80",x"9C",x"45",x"26",x"F8",x"9E",x"41",x"9F", -- 0x2CE0
    x"1B",x"8D",x"36",x"8D",x"02",x"20",x"8D",x"9E", -- 0x2CE8
    x"19",x"EC",x"84",x"27",x"21",x"33",x"04",x"A6", -- 0x2CF0
    x"C0",x"26",x"FC",x"EF",x"84",x"AE",x"84",x"20", -- 0x2CF8
    x"F0",x"DC",x"2B",x"9E",x"19",x"EE",x"84",x"27", -- 0x2D00
    x"09",x"10",x"A3",x"02",x"23",x"06",x"AE",x"84", -- 0x2D08
    x"20",x"F3",x"1A",x"01",x"9F",x"47",x"39",x"26", -- 0x2D10
    x"FB",x"9E",x"19",x"6F",x"80",x"6F",x"80",x"9F", -- 0x2D18
    x"1B",x"9E",x"19",x"BD",x"AE",x"BB",x"9E",x"27", -- 0x2D20
    x"9F",x"23",x"BD",x"AD",x"E4",x"9E",x"1B",x"9F", -- 0x2D28
    x"1D",x"9F",x"1F",x"8E",x"01",x"A9",x"9F",x"0B", -- 0x2D30
    x"AE",x"E4",x"10",x"DE",x"21",x"6F",x"E2",x"0F", -- 0x2D38
    x"2D",x"0F",x"2E",x"0F",x"08",x"6E",x"84",x"86", -- 0x2D40
    x"80",x"97",x"08",x"BD",x"AF",x"89",x"BD",x"AB", -- 0x2D48
    x"F9",x"32",x"62",x"26",x"04",x"9E",x"0F",x"32", -- 0x2D50
    x"85",x"C6",x"09",x"BD",x"AC",x"33",x"BD",x"AE", -- 0x2D58
    x"E8",x"DC",x"68",x"34",x"16",x"C6",x"A5",x"BD", -- 0x2D60
    x"B2",x"6F",x"BD",x"B1",x"43",x"BD",x"B1",x"41", -- 0x2D68
    x"D6",x"54",x"CA",x"7F",x"D4",x"50",x"D7",x"50", -- 0x2D70
    x"10",x"8E",x"AD",x"7F",x"7E",x"B1",x"EA",x"8E", -- 0x2D78
    x"BA",x"C5",x"BD",x"BC",x"14",x"9D",x"A5",x"81", -- 0x2D80
    x"A9",x"26",x"05",x"9D",x"9F",x"BD",x"B1",x"41", -- 0x2D88
    x"BD",x"BC",x"6D",x"BD",x"B1",x"E6",x"DC",x"3B", -- 0x2D90
    x"34",x"06",x"86",x"80",x"34",x"02",x"BD",x"01", -- 0x2D98
    x"9A",x"1C",x"AF",x"8D",x"46",x"9E",x"A6",x"9F", -- 0x2DA0
    x"2F",x"A6",x"80",x"27",x"07",x"81",x"3A",x"27", -- 0x2DA8
    x"0F",x"7E",x"B2",x"77",x"A6",x"81",x"97",x"00", -- 0x2DB0
    x"27",x"5B",x"EC",x"80",x"DD",x"68",x"9F",x"A6", -- 0x2DB8
    x"9D",x"9F",x"8D",x"02",x"20",x"D8",x"27",x"78", -- 0x2DC0
    x"4D",x"10",x"2A",x"01",x"BC",x"81",x"A3",x"22", -- 0x2DC8
    x"0B",x"BE",x"01",x"23",x"48",x"1F",x"89",x"3A", -- 0x2DD0
    x"9D",x"9F",x"6E",x"94",x"81",x"B4",x"23",x"D1", -- 0x2DD8
    x"6E",x"9F",x"01",x"2D",x"9E",x"19",x"30",x"1F", -- 0x2DE0
    x"9F",x"33",x"39",x"BD",x"A1",x"C1",x"27",x"0A", -- 0x2DE8
    x"81",x"03",x"27",x"15",x"81",x"13",x"27",x"03", -- 0x2DF0
    x"97",x"87",x"39",x"BD",x"A1",x"CB",x"27",x"FB", -- 0x2DF8
    x"20",x"EE",x"BD",x"A4",x"26",x"9D",x"A5",x"20", -- 0x2E00
    x"02",x"1A",x"01",x"26",x"33",x"9E",x"A6",x"9F", -- 0x2E08
    x"2F",x"06",x"00",x"32",x"62",x"9E",x"68",x"8C", -- 0x2E10
    x"FF",x"FF",x"27",x"06",x"9F",x"29",x"9E",x"2F", -- 0x2E18
    x"9F",x"2D",x"0F",x"6F",x"8E",x"AB",x"F1",x"0D", -- 0x2E20
    x"00",x"10",x"2A",x"FE",x"46",x"7E",x"AC",x"68", -- 0x2E28
    x"26",x"0E",x"C6",x"20",x"9E",x"2D",x"10",x"27", -- 0x2E30
    x"FE",x"0C",x"9F",x"A6",x"9E",x"29",x"9F",x"68", -- 0x2E38
    x"39",x"27",x"2C",x"BD",x"B3",x"E6",x"34",x"06", -- 0x2E40
    x"9E",x"27",x"9D",x"A5",x"27",x"0C",x"BD",x"B2", -- 0x2E48
    x"6D",x"BD",x"B7",x"3D",x"30",x"1F",x"9C",x"74", -- 0x2E50
    x"22",x"18",x"1F",x"10",x"A3",x"E1",x"25",x"12", -- 0x2E58
    x"1F",x"03",x"83",x"00",x"3A",x"25",x"0B",x"93", -- 0x2E60
    x"1B",x"25",x"07",x"DF",x"21",x"9F",x"27",x"7E", -- 0x2E68
    x"AD",x"26",x"7E",x"AC",x"44",x"BD",x"01",x"94", -- 0x2E70
    x"BD",x"A4",x"26",x"9D",x"A5",x"10",x"27",x"FE", -- 0x2E78
    x"A0",x"BD",x"AD",x"26",x"20",x"19",x"1F",x"89", -- 0x2E80
    x"9D",x"9F",x"C1",x"A5",x"27",x"16",x"C1",x"A6", -- 0x2E88
    x"26",x"45",x"C6",x"03",x"BD",x"AC",x"33",x"DE", -- 0x2E90
    x"A6",x"9E",x"68",x"86",x"A6",x"34",x"52",x"8D", -- 0x2E98
    x"03",x"7E",x"AD",x"9E",x"9D",x"A5",x"BD",x"AF", -- 0x2EA0
    x"67",x"8D",x"40",x"30",x"01",x"DC",x"2B",x"10", -- 0x2EA8
    x"93",x"68",x"22",x"02",x"9E",x"19",x"BD",x"AD", -- 0x2EB0
    x"05",x"25",x"17",x"30",x"1F",x"9F",x"A6",x"39", -- 0x2EB8
    x"26",x"FD",x"86",x"FF",x"97",x"3B",x"BD",x"AB", -- 0x2EC0
    x"F9",x"1F",x"14",x"81",x"26",x"27",x"0B",x"C6", -- 0x2EC8
    x"04",x"8C",x"C6",x"0E",x"7E",x"AC",x"46",x"7E", -- 0x2ED0
    x"B2",x"77",x"35",x"52",x"9F",x"68",x"DF",x"A6", -- 0x2ED8
    x"8D",x"06",x"8C",x"8D",x"06",x"9F",x"A6",x"39", -- 0x2EE0
    x"C6",x"3A",x"86",x"5F",x"D7",x"01",x"5F",x"9E", -- 0x2EE8
    x"A6",x"1F",x"98",x"D6",x"01",x"97",x"01",x"A6", -- 0x2EF0
    x"84",x"27",x"EC",x"34",x"04",x"A1",x"E0",x"27", -- 0x2EF8
    x"E6",x"30",x"01",x"81",x"22",x"27",x"EA",x"4C", -- 0x2F00
    x"26",x"02",x"30",x"01",x"81",x"86",x"26",x"E7", -- 0x2F08
    x"0C",x"04",x"20",x"E3",x"BD",x"B1",x"41",x"9D", -- 0x2F10
    x"A5",x"81",x"81",x"27",x"05",x"C6",x"A7",x"BD", -- 0x2F18
    x"B2",x"6F",x"96",x"4F",x"26",x"13",x"0F",x"04", -- 0x2F20
    x"8D",x"B6",x"4D",x"27",x"BA",x"9D",x"9F",x"81", -- 0x2F28
    x"84",x"26",x"F5",x"0A",x"04",x"2A",x"F1",x"9D", -- 0x2F30
    x"9F",x"9D",x"A5",x"10",x"25",x"FF",x"65",x"7E", -- 0x2F38
    x"AD",x"C6",x"BD",x"B7",x"0B",x"C6",x"81",x"BD", -- 0x2F40
    x"B2",x"6F",x"34",x"02",x"81",x"A6",x"27",x"04", -- 0x2F48
    x"81",x"A5",x"26",x"83",x"0A",x"53",x"26",x"05", -- 0x2F50
    x"35",x"04",x"7E",x"AE",x"88",x"9D",x"9F",x"8D", -- 0x2F58
    x"06",x"81",x"2C",x"27",x"EF",x"35",x"84",x"9E", -- 0x2F60
    x"8A",x"9F",x"2B",x"24",x"61",x"80",x"30",x"97", -- 0x2F68
    x"01",x"DC",x"2B",x"81",x"18",x"22",x"DB",x"58", -- 0x2F70
    x"49",x"58",x"49",x"D3",x"2B",x"58",x"49",x"DB", -- 0x2F78
    x"01",x"89",x"00",x"DD",x"2B",x"9D",x"9F",x"20", -- 0x2F80
    x"E2",x"BD",x"B3",x"57",x"9F",x"3B",x"C6",x"B3", -- 0x2F88
    x"BD",x"B2",x"6F",x"96",x"06",x"34",x"02",x"BD", -- 0x2F90
    x"B1",x"56",x"35",x"02",x"46",x"BD",x"B1",x"48", -- 0x2F98
    x"10",x"27",x"0C",x"8F",x"9E",x"52",x"DC",x"21", -- 0x2FA0
    x"10",x"A3",x"02",x"24",x"11",x"9C",x"1B",x"25", -- 0x2FA8
    x"0D",x"E6",x"84",x"BD",x"B5",x"0D",x"9E",x"4D", -- 0x2FB0
    x"BD",x"B6",x"43",x"8E",x"00",x"56",x"9F",x"4D", -- 0x2FB8
    x"BD",x"B6",x"75",x"DE",x"4D",x"9E",x"3B",x"37", -- 0x2FC0
    x"26",x"A7",x"84",x"10",x"AF",x"02",x"39",x"3F", -- 0x2FC8
    x"52",x"45",x"44",x"4F",x"0D",x"00",x"C6",x"22", -- 0x2FD0
    x"0D",x"6F",x"27",x"03",x"7E",x"AC",x"46",x"96", -- 0x2FD8
    x"09",x"27",x"07",x"9E",x"31",x"9F",x"68",x"7E", -- 0x2FE0
    x"B2",x"77",x"8E",x"AF",x"CE",x"BD",x"B9",x"9C", -- 0x2FE8
    x"9E",x"2F",x"9F",x"A6",x"39",x"C6",x"16",x"9E", -- 0x2FF0
    x"68",x"30",x"01",x"27",x"DF",x"8D",x"03",x"0F", -- 0x2FF8
    x"6F",x"39",x"81",x"23",x"26",x"09",x"BD",x"A5", -- 0x3000
    x"A5",x"BD",x"A3",x"ED",x"BD",x"B2",x"6D",x"81", -- 0x3008
    x"22",x"26",x"0B",x"BD",x"B2",x"44",x"C6",x"3B", -- 0x3010
    x"BD",x"B2",x"6F",x"BD",x"B9",x"9F",x"8E",x"02", -- 0x3018
    x"DC",x"6F",x"84",x"0D",x"6F",x"26",x"22",x"8D", -- 0x3020
    x"06",x"C6",x"2C",x"E7",x"84",x"20",x"1A",x"BD", -- 0x3028
    x"B9",x"AF",x"BD",x"B9",x"AC",x"BD",x"A3",x"90", -- 0x3030
    x"24",x"05",x"32",x"64",x"7E",x"AE",x"11",x"C6", -- 0x3038
    x"2E",x"0D",x"70",x"26",x"97",x"39",x"9E",x"33", -- 0x3040
    x"86",x"4F",x"97",x"09",x"9F",x"35",x"BD",x"B3", -- 0x3048
    x"57",x"9F",x"3B",x"9E",x"A6",x"9F",x"2B",x"9E", -- 0x3050
    x"35",x"A6",x"84",x"26",x"0C",x"96",x"09",x"26", -- 0x3058
    x"58",x"BD",x"01",x"7C",x"BD",x"B9",x"AF",x"8D", -- 0x3060
    x"C6",x"9F",x"A6",x"9D",x"9F",x"D6",x"06",x"27", -- 0x3068
    x"27",x"9E",x"A6",x"97",x"01",x"81",x"22",x"27", -- 0x3070
    x"12",x"30",x"1F",x"4F",x"97",x"01",x"BD",x"A3", -- 0x3078
    x"5F",x"0D",x"6E",x"26",x"06",x"86",x"3A",x"97", -- 0x3080
    x"01",x"86",x"2C",x"97",x"02",x"BD",x"B5",x"1E", -- 0x3088
    x"BD",x"B2",x"49",x"BD",x"AF",x"A4",x"20",x"06", -- 0x3090
    x"BD",x"BD",x"12",x"BD",x"BC",x"33",x"9D",x"A5", -- 0x3098
    x"27",x"06",x"81",x"2C",x"10",x"26",x"FF",x"2E", -- 0x30A0
    x"9E",x"A6",x"9F",x"35",x"9E",x"2B",x"9F",x"A6", -- 0x30A8
    x"9D",x"A5",x"27",x"21",x"BD",x"B2",x"6D",x"20", -- 0x30B0
    x"95",x"9F",x"A6",x"BD",x"AE",x"E8",x"30",x"01", -- 0x30B8
    x"4D",x"26",x"0A",x"C6",x"06",x"EE",x"81",x"27", -- 0x30C0
    x"41",x"EC",x"81",x"DD",x"31",x"A6",x"84",x"81", -- 0x30C8
    x"86",x"26",x"E6",x"20",x"94",x"9E",x"35",x"D6", -- 0x30D0
    x"09",x"10",x"26",x"FD",x"0B",x"A6",x"84",x"27", -- 0x30D8
    x"06",x"8E",x"B0",x"E7",x"7E",x"B9",x"9C",x"39", -- 0x30E0
    x"3F",x"45",x"58",x"54",x"52",x"41",x"20",x"49", -- 0x30E8
    x"47",x"4E",x"4F",x"52",x"45",x"44",x"0D",x"00", -- 0x30F0
    x"26",x"04",x"9E",x"8A",x"20",x"03",x"BD",x"B3", -- 0x30F8
    x"57",x"9F",x"3B",x"BD",x"AB",x"F9",x"27",x"04", -- 0x3100
    x"C6",x"00",x"20",x"47",x"1F",x"14",x"30",x"03", -- 0x3108
    x"BD",x"BC",x"14",x"A6",x"68",x"97",x"54",x"9E", -- 0x3110
    x"3B",x"BD",x"B9",x"C2",x"BD",x"BC",x"33",x"30", -- 0x3118
    x"69",x"BD",x"BC",x"96",x"E0",x"68",x"27",x"0C", -- 0x3120
    x"AE",x"6E",x"9F",x"68",x"AE",x"E8",x"10",x"9F", -- 0x3128
    x"A6",x"7E",x"AD",x"9E",x"32",x"E8",x"12",x"9D", -- 0x3130
    x"A5",x"81",x"2C",x"26",x"F4",x"9D",x"9F",x"8D", -- 0x3138
    x"BD",x"8D",x"13",x"1C",x"FE",x"7D",x"1A",x"01", -- 0x3140
    x"0D",x"06",x"25",x"03",x"2A",x"99",x"8C",x"2B", -- 0x3148
    x"96",x"C6",x"18",x"7E",x"AC",x"46",x"8D",x"6E", -- 0x3150
    x"4F",x"8C",x"34",x"04",x"34",x"02",x"C6",x"01", -- 0x3158
    x"BD",x"AC",x"33",x"BD",x"B2",x"23",x"0F",x"3F", -- 0x3160
    x"9D",x"A5",x"80",x"B2",x"25",x"13",x"81",x"03", -- 0x3168
    x"24",x"0F",x"81",x"01",x"49",x"98",x"3F",x"91", -- 0x3170
    x"3F",x"25",x"64",x"97",x"3F",x"9D",x"9F",x"20", -- 0x3178
    x"E9",x"D6",x"3F",x"26",x"33",x"10",x"24",x"00", -- 0x3180
    x"6B",x"8B",x"07",x"24",x"67",x"99",x"06",x"10", -- 0x3188
    x"27",x"04",x"7C",x"89",x"FF",x"34",x"02",x"48", -- 0x3190
    x"AB",x"E0",x"8E",x"AA",x"51",x"30",x"86",x"35", -- 0x3198
    x"02",x"A1",x"84",x"24",x"55",x"8D",x"9C",x"34", -- 0x31A0
    x"02",x"8D",x"29",x"9E",x"3D",x"35",x"02",x"26", -- 0x31A8
    x"1D",x"4D",x"10",x"27",x"00",x"6A",x"20",x"4B", -- 0x31B0
    x"08",x"06",x"59",x"8D",x"09",x"8E",x"B1",x"CB", -- 0x31B8
    x"D7",x"3F",x"0F",x"06",x"20",x"D9",x"9E",x"A6", -- 0x31C0
    x"7E",x"AE",x"BB",x"64",x"B2",x"F4",x"A1",x"84", -- 0x31C8
    x"24",x"31",x"20",x"D3",x"EC",x"01",x"34",x"06", -- 0x31D0
    x"8D",x"08",x"D6",x"3F",x"16",x"FF",x"7B",x"7E", -- 0x31D8
    x"B2",x"77",x"D6",x"54",x"A6",x"84",x"35",x"20", -- 0x31E0
    x"34",x"04",x"D6",x"4F",x"9E",x"50",x"DE",x"52", -- 0x31E8
    x"34",x"54",x"6E",x"A4",x"9E",x"8A",x"A6",x"E0", -- 0x31F0
    x"27",x"26",x"81",x"64",x"27",x"03",x"BD",x"B1", -- 0x31F8
    x"43",x"9F",x"3D",x"35",x"04",x"81",x"5A",x"27", -- 0x3200
    x"19",x"81",x"7D",x"27",x"15",x"54",x"D7",x"0A", -- 0x3208
    x"35",x"52",x"97",x"5C",x"9F",x"5D",x"DF",x"5F", -- 0x3210
    x"35",x"04",x"D7",x"61",x"D8",x"54",x"D7",x"62", -- 0x3218
    x"D6",x"4F",x"39",x"BD",x"01",x"8B",x"0F",x"06", -- 0x3220
    x"9D",x"9F",x"24",x"03",x"7E",x"BD",x"12",x"BD", -- 0x3228
    x"B3",x"A2",x"24",x"50",x"81",x"2E",x"27",x"F4", -- 0x3230
    x"81",x"AC",x"27",x"40",x"81",x"AB",x"27",x"E3", -- 0x3238
    x"81",x"22",x"26",x"0A",x"9E",x"A6",x"BD",x"B5", -- 0x3240
    x"18",x"9E",x"64",x"9F",x"A6",x"39",x"81",x"A8", -- 0x3248
    x"26",x"0D",x"86",x"5A",x"BD",x"B1",x"5A",x"BD", -- 0x3250
    x"B3",x"ED",x"43",x"53",x"7E",x"B4",x"F4",x"4C", -- 0x3258
    x"27",x"2E",x"8D",x"06",x"BD",x"B1",x"56",x"C6", -- 0x3260
    x"29",x"8C",x"C6",x"28",x"8C",x"C6",x"2C",x"E1", -- 0x3268
    x"9F",x"00",x"A6",x"26",x"02",x"0E",x"9F",x"C6", -- 0x3270
    x"02",x"7E",x"AC",x"46",x"86",x"7D",x"BD",x"B1", -- 0x3278
    x"5A",x"7E",x"BE",x"E9",x"BD",x"B3",x"57",x"9F", -- 0x3280
    x"52",x"96",x"06",x"26",x"95",x"7E",x"BC",x"14", -- 0x3288
    x"9D",x"9F",x"1F",x"89",x"58",x"9D",x"9F",x"C1", -- 0x3290
    x"26",x"23",x"04",x"6E",x"9F",x"01",x"32",x"34", -- 0x3298
    x"04",x"C1",x"1C",x"25",x"22",x"C1",x"24",x"24", -- 0x32A0
    x"20",x"8D",x"BF",x"A6",x"E4",x"81",x"22",x"24", -- 0x32A8
    x"18",x"BD",x"B1",x"56",x"8D",x"B7",x"BD",x"B1", -- 0x32B0
    x"46",x"35",x"02",x"DE",x"52",x"34",x"42",x"BD", -- 0x32B8
    x"B7",x"0B",x"35",x"02",x"34",x"06",x"8E",x"8D", -- 0x32C0
    x"99",x"35",x"04",x"BE",x"01",x"28",x"3A",x"AD", -- 0x32C8
    x"94",x"7E",x"B1",x"43",x"86",x"4F",x"97",x"03", -- 0x32D0
    x"BD",x"B3",x"ED",x"DD",x"01",x"BD",x"BC",x"4A", -- 0x32D8
    x"BD",x"B3",x"ED",x"0D",x"03",x"26",x"06",x"94", -- 0x32E0
    x"01",x"D4",x"02",x"20",x"04",x"9A",x"01",x"DA", -- 0x32E8
    x"02",x"7E",x"B4",x"F4",x"BD",x"B1",x"48",x"26", -- 0x32F0
    x"10",x"96",x"61",x"8A",x"7F",x"94",x"5D",x"97", -- 0x32F8
    x"5D",x"8E",x"00",x"5C",x"BD",x"BC",x"96",x"20", -- 0x3300
    x"36",x"0F",x"06",x"0A",x"3F",x"BD",x"B6",x"57", -- 0x3308
    x"D7",x"56",x"9F",x"58",x"9E",x"5F",x"BD",x"B6", -- 0x3310
    x"59",x"96",x"56",x"34",x"04",x"A0",x"E0",x"27", -- 0x3318
    x"07",x"86",x"01",x"24",x"03",x"D6",x"56",x"40", -- 0x3320
    x"97",x"54",x"DE",x"58",x"5C",x"5A",x"26",x"04", -- 0x3328
    x"D6",x"54",x"20",x"0B",x"A6",x"80",x"A1",x"C0", -- 0x3330
    x"27",x"F3",x"C6",x"FF",x"24",x"01",x"50",x"CB", -- 0x3338
    x"01",x"59",x"D4",x"0A",x"27",x"02",x"C6",x"FF", -- 0x3340
    x"7E",x"BC",x"7C",x"BD",x"B2",x"6D",x"C6",x"01", -- 0x3348
    x"8D",x"08",x"9D",x"A5",x"26",x"F5",x"39",x"5F", -- 0x3350
    x"9D",x"A5",x"D7",x"05",x"97",x"37",x"9D",x"A5", -- 0x3358
    x"8D",x"40",x"10",x"25",x"FF",x"11",x"5F",x"D7", -- 0x3360
    x"06",x"9D",x"9F",x"25",x"04",x"8D",x"33",x"25", -- 0x3368
    x"0A",x"1F",x"89",x"9D",x"9F",x"25",x"FC",x"8D", -- 0x3370
    x"29",x"24",x"F8",x"81",x"24",x"26",x"06",x"03", -- 0x3378
    x"06",x"CB",x"80",x"9D",x"9F",x"D7",x"38",x"9A", -- 0x3380
    x"08",x"80",x"28",x"10",x"27",x"00",x"75",x"0F", -- 0x3388
    x"08",x"9E",x"1B",x"DC",x"37",x"9C",x"1D",x"27", -- 0x3390
    x"12",x"10",x"A3",x"81",x"27",x"3E",x"30",x"05", -- 0x3398
    x"20",x"F3",x"81",x"41",x"25",x"04",x"80",x"5B", -- 0x33A0
    x"80",x"A5",x"39",x"8E",x"00",x"8A",x"EE",x"E4", -- 0x33A8
    x"11",x"83",x"B2",x"87",x"27",x"28",x"DC",x"1F", -- 0x33B0
    x"DD",x"43",x"C3",x"00",x"07",x"DD",x"41",x"9E", -- 0x33B8
    x"1D",x"9F",x"47",x"BD",x"AC",x"1E",x"9E",x"41", -- 0x33C0
    x"9F",x"1F",x"9E",x"45",x"9F",x"1D",x"9E",x"47", -- 0x33C8
    x"DC",x"37",x"ED",x"81",x"4F",x"5F",x"ED",x"84", -- 0x33D0
    x"ED",x"02",x"A7",x"04",x"9F",x"39",x"39",x"90", -- 0x33D8
    x"80",x"00",x"00",x"00",x"9D",x"9F",x"BD",x"B1", -- 0x33E0
    x"41",x"96",x"54",x"2B",x"5D",x"BD",x"B1",x"43", -- 0x33E8
    x"96",x"4F",x"81",x"90",x"25",x"08",x"8E",x"B3", -- 0x33F0
    x"DF",x"BD",x"BC",x"96",x"26",x"4C",x"BD",x"BC", -- 0x33F8
    x"C8",x"DC",x"52",x"39",x"DC",x"05",x"34",x"06", -- 0x3400
    x"12",x"5F",x"9E",x"37",x"34",x"14",x"8D",x"D4", -- 0x3408
    x"35",x"34",x"9F",x"37",x"DE",x"52",x"34",x"60", -- 0x3410
    x"5C",x"9D",x"A5",x"81",x"2C",x"27",x"EB",x"D7", -- 0x3418
    x"03",x"BD",x"B2",x"67",x"35",x"06",x"DD",x"05", -- 0x3420
    x"9E",x"1D",x"9C",x"1F",x"27",x"21",x"DC",x"37", -- 0x3428
    x"10",x"A3",x"84",x"27",x"06",x"EC",x"02",x"30", -- 0x3430
    x"8B",x"20",x"EF",x"C6",x"12",x"96",x"05",x"26", -- 0x3438
    x"0B",x"D6",x"03",x"E1",x"04",x"27",x"59",x"C6", -- 0x3440
    x"10",x"8C",x"C6",x"08",x"7E",x"AC",x"46",x"CC", -- 0x3448
    x"00",x"05",x"DD",x"64",x"DC",x"37",x"ED",x"84", -- 0x3450
    x"D6",x"03",x"E7",x"04",x"BD",x"AC",x"33",x"9F", -- 0x3458
    x"41",x"C6",x"0B",x"4F",x"0D",x"05",x"27",x"05", -- 0x3460
    x"35",x"06",x"C3",x"00",x"01",x"ED",x"05",x"8D", -- 0x3468
    x"5D",x"DD",x"64",x"30",x"02",x"0A",x"03",x"26", -- 0x3470
    x"E8",x"9F",x"0F",x"D3",x"0F",x"10",x"25",x"F7", -- 0x3478
    x"C3",x"1F",x"01",x"BD",x"AC",x"37",x"83",x"00", -- 0x3480
    x"35",x"DD",x"1F",x"4F",x"30",x"1F",x"A7",x"05", -- 0x3488
    x"9C",x"0F",x"26",x"F8",x"9E",x"41",x"96",x"1F", -- 0x3490
    x"93",x"41",x"ED",x"02",x"96",x"05",x"26",x"2D", -- 0x3498
    x"E6",x"04",x"D7",x"03",x"4F",x"5F",x"DD",x"64", -- 0x34A0
    x"35",x"06",x"DD",x"52",x"10",x"A3",x"05",x"24", -- 0x34A8
    x"3A",x"DE",x"64",x"27",x"04",x"8D",x"17",x"D3", -- 0x34B0
    x"52",x"30",x"02",x"0A",x"03",x"26",x"E7",x"ED", -- 0x34B8
    x"E3",x"58",x"49",x"58",x"49",x"E3",x"E1",x"30", -- 0x34C0
    x"8B",x"30",x"05",x"9F",x"39",x"39",x"86",x"10", -- 0x34C8
    x"97",x"45",x"EC",x"05",x"DD",x"17",x"4F",x"5F", -- 0x34D0
    x"58",x"49",x"25",x"0F",x"08",x"65",x"09",x"64", -- 0x34D8
    x"24",x"04",x"D3",x"17",x"25",x"05",x"0A",x"45", -- 0x34E0
    x"26",x"EE",x"39",x"7E",x"B4",x"47",x"1F",x"40", -- 0x34E8
    x"93",x"1F",x"21",x"4F",x"0F",x"06",x"DD",x"50", -- 0x34F0
    x"C6",x"90",x"7E",x"BC",x"82",x"BD",x"B1",x"43", -- 0x34F8
    x"CE",x"03",x"D9",x"BD",x"BD",x"DC",x"32",x"62", -- 0x3500
    x"8E",x"03",x"D8",x"20",x"0B",x"9F",x"4D",x"8D", -- 0x3508
    x"5C",x"9F",x"58",x"D7",x"56",x"39",x"30",x"1F", -- 0x3510
    x"86",x"22",x"97",x"01",x"97",x"02",x"30",x"01", -- 0x3518
    x"9F",x"62",x"9F",x"58",x"C6",x"FF",x"5C",x"A6", -- 0x3520
    x"80",x"27",x"0C",x"91",x"01",x"27",x"04",x"91", -- 0x3528
    x"02",x"26",x"F3",x"81",x"22",x"27",x"02",x"30", -- 0x3530
    x"1F",x"9F",x"64",x"D7",x"56",x"DE",x"62",x"11", -- 0x3538
    x"83",x"03",x"D9",x"22",x"07",x"8D",x"C6",x"9E", -- 0x3540
    x"62",x"BD",x"B6",x"45",x"9E",x"0B",x"8C",x"01", -- 0x3548
    x"D1",x"26",x"05",x"C6",x"1E",x"7E",x"AC",x"46", -- 0x3550
    x"96",x"56",x"A7",x"00",x"DC",x"58",x"ED",x"02", -- 0x3558
    x"86",x"FF",x"97",x"06",x"9F",x"0D",x"9F",x"52", -- 0x3560
    x"30",x"05",x"9F",x"0B",x"39",x"0F",x"07",x"4F", -- 0x3568
    x"34",x"06",x"DC",x"23",x"A3",x"E0",x"10",x"93", -- 0x3570
    x"21",x"25",x"0A",x"DD",x"23",x"9E",x"23",x"30", -- 0x3578
    x"01",x"9F",x"25",x"35",x"84",x"C6",x"1A",x"03", -- 0x3580
    x"07",x"27",x"CA",x"8D",x"04",x"35",x"04",x"20", -- 0x3588
    x"DE",x"9E",x"27",x"9F",x"23",x"4F",x"5F",x"DD", -- 0x3590
    x"4B",x"9E",x"21",x"9F",x"47",x"8E",x"01",x"A9", -- 0x3598
    x"9C",x"0B",x"27",x"04",x"8D",x"32",x"20",x"F8", -- 0x35A0
    x"9E",x"1B",x"9C",x"1D",x"27",x"04",x"8D",x"22", -- 0x35A8
    x"20",x"F8",x"9F",x"41",x"9E",x"41",x"9C",x"1F", -- 0x35B0
    x"27",x"35",x"EC",x"02",x"D3",x"41",x"DD",x"41", -- 0x35B8
    x"A6",x"01",x"2A",x"F0",x"E6",x"04",x"58",x"CB", -- 0x35C0
    x"05",x"3A",x"9C",x"41",x"27",x"E8",x"8D",x"08", -- 0x35C8
    x"20",x"F8",x"A6",x"01",x"30",x"02",x"2A",x"14", -- 0x35D0
    x"E6",x"84",x"27",x"10",x"EC",x"02",x"10",x"93", -- 0x35D8
    x"23",x"22",x"09",x"10",x"93",x"47",x"23",x"04", -- 0x35E0
    x"9F",x"4B",x"DD",x"47",x"30",x"05",x"39",x"9E", -- 0x35E8
    x"4B",x"27",x"FB",x"4F",x"E6",x"84",x"5A",x"D3", -- 0x35F0
    x"47",x"DD",x"43",x"9E",x"23",x"9F",x"41",x"BD", -- 0x35F8
    x"AC",x"20",x"9E",x"4B",x"DC",x"45",x"ED",x"02", -- 0x3600
    x"9E",x"45",x"30",x"1F",x"7E",x"B5",x"93",x"DC", -- 0x3608
    x"52",x"34",x"06",x"BD",x"B2",x"23",x"BD",x"B1", -- 0x3610
    x"46",x"35",x"10",x"9F",x"62",x"E6",x"84",x"9E", -- 0x3618
    x"52",x"EB",x"84",x"24",x"05",x"C6",x"1C",x"7E", -- 0x3620
    x"AC",x"46",x"BD",x"B5",x"0D",x"9E",x"62",x"E6", -- 0x3628
    x"84",x"8D",x"10",x"9E",x"4D",x"8D",x"22",x"8D", -- 0x3630
    x"0C",x"9E",x"62",x"8D",x"1C",x"BD",x"B5",x"4C", -- 0x3638
    x"7E",x"B1",x"68",x"AE",x"02",x"DE",x"25",x"5C", -- 0x3640
    x"20",x"04",x"A6",x"80",x"A7",x"C0",x"5A",x"26", -- 0x3648
    x"F9",x"DF",x"25",x"39",x"BD",x"B1",x"46",x"9E", -- 0x3650
    x"52",x"E6",x"84",x"8D",x"18",x"26",x"13",x"AE", -- 0x3658
    x"07",x"30",x"1F",x"9C",x"23",x"26",x"08",x"34", -- 0x3660
    x"04",x"D3",x"23",x"DD",x"23",x"35",x"04",x"30", -- 0x3668
    x"01",x"39",x"AE",x"02",x"39",x"9C",x"0D",x"26", -- 0x3670
    x"07",x"9F",x"0B",x"30",x"1B",x"9F",x"0D",x"4F", -- 0x3678
    x"39",x"8D",x"03",x"7E",x"B4",x"F3",x"8D",x"CC", -- 0x3680
    x"0F",x"06",x"5D",x"39",x"BD",x"B7",x"0E",x"C6", -- 0x3688
    x"01",x"BD",x"B5",x"6D",x"96",x"53",x"BD",x"B5", -- 0x3690
    x"11",x"A7",x"84",x"32",x"62",x"7E",x"B5",x"4C", -- 0x3698
    x"8D",x"02",x"20",x"DF",x"8D",x"E0",x"27",x"5E", -- 0x36A0
    x"E6",x"84",x"39",x"8D",x"48",x"4F",x"E1",x"84", -- 0x36A8
    x"23",x"03",x"E6",x"84",x"4F",x"34",x"06",x"BD", -- 0x36B0
    x"B5",x"0F",x"9E",x"4D",x"8D",x"9B",x"35",x"04", -- 0x36B8
    x"3A",x"35",x"04",x"BD",x"B6",x"45",x"20",x"D5", -- 0x36C0
    x"8D",x"2B",x"A0",x"84",x"40",x"20",x"DF",x"C6", -- 0x36C8
    x"FF",x"D7",x"53",x"9D",x"A5",x"81",x"29",x"27", -- 0x36D0
    x"05",x"BD",x"B2",x"6D",x"8D",x"2D",x"8D",x"15", -- 0x36D8
    x"27",x"24",x"5F",x"4A",x"A1",x"84",x"24",x"CD", -- 0x36E0
    x"1F",x"89",x"E0",x"84",x"50",x"D1",x"53",x"23", -- 0x36E8
    x"C4",x"D6",x"53",x"20",x"C0",x"BD",x"B2",x"67", -- 0x36F0
    x"EE",x"E4",x"AE",x"65",x"9F",x"4D",x"A6",x"64", -- 0x36F8
    x"E6",x"64",x"32",x"67",x"1F",x"35",x"7E",x"B4", -- 0x3700
    x"4A",x"9D",x"9F",x"BD",x"B1",x"41",x"BD",x"B3", -- 0x3708
    x"E9",x"4D",x"26",x"F2",x"0E",x"A5",x"BD",x"B6", -- 0x3710
    x"86",x"10",x"27",x"03",x"1C",x"DE",x"A6",x"9F", -- 0x3718
    x"A6",x"3A",x"A6",x"84",x"34",x"52",x"6F",x"84", -- 0x3720
    x"9D",x"A5",x"BD",x"BD",x"12",x"35",x"52",x"A7", -- 0x3728
    x"84",x"DF",x"A6",x"39",x"8D",x"07",x"9F",x"2B", -- 0x3730
    x"BD",x"B2",x"6D",x"20",x"CE",x"BD",x"B1",x"41", -- 0x3738
    x"96",x"54",x"2B",x"C2",x"96",x"4F",x"81",x"90", -- 0x3740
    x"22",x"BC",x"BD",x"BC",x"C8",x"9E",x"52",x"39", -- 0x3748
    x"8D",x"EE",x"E6",x"84",x"7E",x"B4",x"F3",x"8D", -- 0x3750
    x"DB",x"9E",x"2B",x"E7",x"84",x"39",x"C6",x"FE", -- 0x3758
    x"D7",x"6F",x"9D",x"A5",x"34",x"01",x"BD",x"AF", -- 0x3760
    x"67",x"BD",x"AD",x"01",x"9F",x"66",x"35",x"01", -- 0x3768
    x"27",x"12",x"9D",x"A5",x"27",x"13",x"81",x"AC", -- 0x3770
    x"26",x"09",x"9D",x"9F",x"27",x"06",x"BD",x"AF", -- 0x3778
    x"67",x"27",x"06",x"39",x"CE",x"FF",x"FF",x"DF", -- 0x3780
    x"2B",x"32",x"62",x"9E",x"66",x"BD",x"B9",x"5C", -- 0x3788
    x"BD",x"A5",x"49",x"EC",x"84",x"26",x"08",x"BD", -- 0x3790
    x"A4",x"2D",x"0F",x"6F",x"7E",x"AC",x"73",x"9F", -- 0x3798
    x"66",x"EC",x"02",x"10",x"93",x"2B",x"22",x"EF", -- 0x37A0
    x"BD",x"BD",x"CC",x"BD",x"B9",x"AC",x"9E",x"66", -- 0x37A8
    x"8D",x"10",x"AE",x"9F",x"00",x"66",x"CE",x"02", -- 0x37B0
    x"DD",x"A6",x"C0",x"27",x"D0",x"BD",x"B9",x"B1", -- 0x37B8
    x"20",x"F7",x"BD",x"01",x"A6",x"30",x"04",x"10", -- 0x37C0
    x"8E",x"02",x"DD",x"A6",x"80",x"27",x"51",x"2B", -- 0x37C8
    x"15",x"81",x"3A",x"26",x"0D",x"E6",x"84",x"C1", -- 0x37D0
    x"84",x"27",x"F0",x"C1",x"83",x"27",x"EC",x"8C", -- 0x37D8
    x"86",x"21",x"8D",x"30",x"20",x"E5",x"CE",x"01", -- 0x37E0
    x"16",x"81",x"FF",x"26",x"04",x"A6",x"80",x"33", -- 0x37E8
    x"45",x"84",x"7F",x"33",x"4A",x"6D",x"C4",x"27", -- 0x37F0
    x"E7",x"A0",x"C4",x"2A",x"F6",x"AB",x"C4",x"EE", -- 0x37F8
    x"41",x"4A",x"2B",x"06",x"6D",x"C0",x"2A",x"FC", -- 0x3800
    x"20",x"F7",x"A6",x"C4",x"8D",x"06",x"6D",x"C0", -- 0x3808
    x"2A",x"F8",x"20",x"B7",x"10",x"8C",x"03",x"D6", -- 0x3810
    x"24",x"06",x"84",x"7F",x"A7",x"A0",x"6F",x"A4", -- 0x3818
    x"39",x"BD",x"01",x"A3",x"9E",x"A6",x"CE",x"02", -- 0x3820
    x"DC",x"0F",x"43",x"0F",x"44",x"A6",x"80",x"27", -- 0x3828
    x"21",x"0D",x"43",x"27",x"0F",x"BD",x"B3",x"A2", -- 0x3830
    x"24",x"18",x"81",x"30",x"25",x"04",x"81",x"39", -- 0x3838
    x"23",x"10",x"0F",x"43",x"81",x"20",x"27",x"0A", -- 0x3840
    x"97",x"42",x"81",x"22",x"27",x"38",x"0D",x"44", -- 0x3848
    x"27",x"19",x"A7",x"C0",x"27",x"06",x"81",x"3A", -- 0x3850
    x"27",x"CF",x"20",x"D1",x"6F",x"C0",x"6F",x"C0", -- 0x3858
    x"1F",x"30",x"83",x"02",x"DA",x"8E",x"02",x"DB", -- 0x3860
    x"9F",x"A6",x"39",x"81",x"3F",x"26",x"04",x"86", -- 0x3868
    x"87",x"20",x"DF",x"81",x"27",x"26",x"13",x"CC", -- 0x3870
    x"3A",x"83",x"ED",x"C1",x"0F",x"42",x"A6",x"80", -- 0x3878
    x"27",x"D0",x"91",x"42",x"27",x"CC",x"A7",x"C0", -- 0x3880
    x"20",x"F4",x"81",x"30",x"25",x"04",x"81",x"3C", -- 0x3888
    x"25",x"C0",x"30",x"1F",x"34",x"50",x"0F",x"41", -- 0x3890
    x"CE",x"01",x"16",x"0F",x"42",x"33",x"4A",x"A6", -- 0x3898
    x"C4",x"27",x"31",x"10",x"AE",x"41",x"AE",x"E4", -- 0x38A0
    x"E6",x"A0",x"E0",x"80",x"27",x"FA",x"C1",x"80", -- 0x38A8
    x"26",x"38",x"32",x"62",x"35",x"40",x"DA",x"42", -- 0x38B0
    x"96",x"41",x"26",x"06",x"C1",x"84",x"26",x"06", -- 0x38B8
    x"86",x"3A",x"ED",x"C1",x"20",x"94",x"E7",x"C0", -- 0x38C0
    x"C1",x"86",x"26",x"02",x"0C",x"44",x"C1",x"82", -- 0x38C8
    x"27",x"AA",x"20",x"86",x"CE",x"01",x"1B",x"03", -- 0x38D0
    x"41",x"26",x"C0",x"35",x"50",x"A6",x"80",x"A7", -- 0x38D8
    x"C0",x"BD",x"B3",x"A2",x"25",x"EC",x"03",x"43", -- 0x38E0
    x"20",x"E8",x"0C",x"42",x"4A",x"27",x"AE",x"31", -- 0x38E8
    x"3F",x"E6",x"A0",x"2A",x"FC",x"20",x"AF",x"27", -- 0x38F0
    x"5F",x"8D",x"03",x"0F",x"6F",x"39",x"81",x"40", -- 0x38F8
    x"26",x"05",x"BD",x"A5",x"54",x"20",x"0A",x"81", -- 0x3900
    x"23",x"26",x"0D",x"BD",x"A5",x"A5",x"BD",x"A4", -- 0x3908
    x"06",x"9D",x"A5",x"27",x"43",x"BD",x"B2",x"6D", -- 0x3910
    x"BD",x"01",x"79",x"27",x"48",x"81",x"A4",x"27", -- 0x3918
    x"5D",x"81",x"2C",x"27",x"41",x"81",x"3B",x"27", -- 0x3920
    x"6E",x"BD",x"B1",x"56",x"96",x"06",x"34",x"02", -- 0x3928
    x"26",x"06",x"BD",x"BD",x"D9",x"BD",x"B5",x"16", -- 0x3930
    x"8D",x"65",x"35",x"04",x"BD",x"A3",x"5F",x"0D", -- 0x3938
    x"6E",x"27",x"06",x"8D",x"13",x"9D",x"A5",x"20", -- 0x3940
    x"D2",x"5D",x"26",x"08",x"9D",x"A5",x"81",x"2C", -- 0x3948
    x"27",x"14",x"8D",x"58",x"9D",x"A5",x"26",x"C5", -- 0x3950
    x"86",x"0D",x"20",x"55",x"BD",x"A3",x"5F",x"27", -- 0x3958
    x"F7",x"96",x"6C",x"26",x"F3",x"39",x"BD",x"A3", -- 0x3960
    x"5F",x"27",x"0A",x"D6",x"6C",x"D1",x"6B",x"25", -- 0x3968
    x"06",x"8D",x"E5",x"20",x"22",x"D6",x"6C",x"D0", -- 0x3970
    x"6A",x"24",x"FC",x"50",x"20",x"10",x"BD",x"B7", -- 0x3978
    x"09",x"81",x"29",x"10",x"26",x"F8",x"F0",x"BD", -- 0x3980
    x"A3",x"5F",x"D0",x"6C",x"23",x"09",x"0D",x"6E", -- 0x3988
    x"26",x"05",x"8D",x"18",x"5A",x"26",x"FB",x"9D", -- 0x3990
    x"9F",x"7E",x"B9",x"1B",x"BD",x"B5",x"18",x"BD", -- 0x3998
    x"B6",x"57",x"5C",x"5A",x"27",x"BF",x"A6",x"80", -- 0x39A0
    x"8D",x"07",x"20",x"F7",x"86",x"20",x"8C",x"86", -- 0x39A8
    x"3F",x"7E",x"A2",x"82",x"8E",x"BE",x"C0",x"20", -- 0x39B0
    x"09",x"BD",x"BB",x"2F",x"03",x"54",x"03",x"62", -- 0x39B8
    x"20",x"03",x"BD",x"BB",x"2F",x"5D",x"10",x"27", -- 0x39C0
    x"02",x"80",x"8E",x"00",x"5C",x"1F",x"89",x"5D", -- 0x39C8
    x"27",x"6C",x"D0",x"4F",x"27",x"69",x"25",x"0A", -- 0x39D0
    x"97",x"4F",x"96",x"61",x"97",x"54",x"8E",x"00", -- 0x39D8
    x"4F",x"50",x"C1",x"F8",x"2F",x"59",x"4F",x"64", -- 0x39E0
    x"01",x"BD",x"BA",x"BA",x"D6",x"62",x"2A",x"0B", -- 0x39E8
    x"63",x"01",x"63",x"02",x"63",x"03",x"63",x"04", -- 0x39F0
    x"43",x"89",x"00",x"97",x"63",x"96",x"53",x"99", -- 0x39F8
    x"60",x"97",x"53",x"96",x"52",x"99",x"5F",x"97", -- 0x3A00
    x"52",x"96",x"51",x"99",x"5E",x"97",x"51",x"96", -- 0x3A08
    x"50",x"99",x"5D",x"97",x"50",x"5D",x"2A",x"44", -- 0x3A10
    x"25",x"02",x"8D",x"5D",x"5F",x"96",x"50",x"26", -- 0x3A18
    x"2E",x"96",x"51",x"97",x"50",x"96",x"52",x"97", -- 0x3A20
    x"51",x"96",x"53",x"97",x"52",x"96",x"63",x"97", -- 0x3A28
    x"53",x"0F",x"63",x"CB",x"08",x"C1",x"28",x"2D", -- 0x3A30
    x"E4",x"4F",x"97",x"4F",x"97",x"54",x"39",x"8D", -- 0x3A38
    x"6D",x"5F",x"20",x"A8",x"5C",x"08",x"63",x"09", -- 0x3A40
    x"53",x"09",x"52",x"09",x"51",x"09",x"50",x"2A", -- 0x3A48
    x"F3",x"96",x"4F",x"34",x"04",x"A0",x"E0",x"97", -- 0x3A50
    x"4F",x"23",x"DE",x"8C",x"25",x"08",x"08",x"63", -- 0x3A58
    x"86",x"00",x"97",x"63",x"20",x"0C",x"0C",x"4F", -- 0x3A60
    x"27",x"28",x"06",x"50",x"06",x"51",x"06",x"52", -- 0x3A68
    x"06",x"53",x"24",x"04",x"8D",x"0D",x"27",x"EE", -- 0x3A70
    x"39",x"03",x"54",x"03",x"50",x"03",x"51",x"03", -- 0x3A78
    x"52",x"03",x"53",x"9E",x"52",x"30",x"01",x"9F", -- 0x3A80
    x"52",x"26",x"06",x"9E",x"50",x"30",x"01",x"9F", -- 0x3A88
    x"50",x"39",x"C6",x"0A",x"7E",x"AC",x"46",x"8E", -- 0x3A90
    x"00",x"12",x"A6",x"04",x"97",x"63",x"A6",x"03", -- 0x3A98
    x"A7",x"04",x"A6",x"02",x"A7",x"03",x"A6",x"01", -- 0x3AA0
    x"A7",x"02",x"96",x"5B",x"A7",x"01",x"CB",x"08", -- 0x3AA8
    x"2F",x"E8",x"96",x"63",x"C0",x"08",x"27",x"0C", -- 0x3AB0
    x"67",x"01",x"66",x"02",x"66",x"03",x"66",x"04", -- 0x3AB8
    x"46",x"5C",x"26",x"F4",x"39",x"81",x"00",x"00", -- 0x3AC0
    x"00",x"00",x"8D",x"63",x"27",x"60",x"8D",x"78", -- 0x3AC8
    x"86",x"00",x"97",x"13",x"97",x"14",x"97",x"15", -- 0x3AD0
    x"97",x"16",x"D6",x"53",x"8D",x"22",x"D6",x"63", -- 0x3AD8
    x"D7",x"AE",x"D6",x"52",x"8D",x"1A",x"D6",x"63", -- 0x3AE0
    x"D7",x"AD",x"D6",x"51",x"8D",x"12",x"D6",x"63", -- 0x3AE8
    x"D7",x"AC",x"D6",x"50",x"8D",x"0C",x"D6",x"63", -- 0x3AF0
    x"D7",x"AB",x"BD",x"BC",x"0B",x"7E",x"BA",x"1C", -- 0x3AF8
    x"27",x"95",x"43",x"96",x"13",x"56",x"27",x"26", -- 0x3B00
    x"24",x"16",x"96",x"16",x"9B",x"60",x"97",x"16", -- 0x3B08
    x"96",x"15",x"99",x"5F",x"97",x"15",x"96",x"14", -- 0x3B10
    x"99",x"5E",x"97",x"14",x"96",x"13",x"99",x"5D", -- 0x3B18
    x"46",x"97",x"13",x"06",x"14",x"06",x"15",x"06", -- 0x3B20
    x"16",x"06",x"63",x"4F",x"20",x"D5",x"39",x"EC", -- 0x3B28
    x"01",x"97",x"61",x"8A",x"80",x"DD",x"5D",x"D6", -- 0x3B30
    x"61",x"D8",x"54",x"D7",x"62",x"EC",x"03",x"DD", -- 0x3B38
    x"5F",x"A6",x"84",x"97",x"5C",x"D6",x"4F",x"39", -- 0x3B40
    x"4D",x"27",x"16",x"9B",x"4F",x"46",x"49",x"28", -- 0x3B48
    x"10",x"8B",x"80",x"97",x"4F",x"27",x"0C",x"96", -- 0x3B50
    x"62",x"97",x"54",x"39",x"96",x"54",x"43",x"20", -- 0x3B58
    x"02",x"32",x"62",x"10",x"2A",x"FE",x"D2",x"7E", -- 0x3B60
    x"BA",x"92",x"BD",x"BC",x"5F",x"27",x"0D",x"8B", -- 0x3B68
    x"02",x"25",x"F4",x"0F",x"62",x"BD",x"B9",x"CD", -- 0x3B70
    x"0C",x"4F",x"27",x"EB",x"39",x"84",x"20",x"00", -- 0x3B78
    x"00",x"00",x"BD",x"BC",x"5F",x"8E",x"BB",x"7D", -- 0x3B80
    x"5F",x"D7",x"62",x"BD",x"BC",x"14",x"8C",x"8D", -- 0x3B88
    x"9E",x"27",x"73",x"00",x"4F",x"8D",x"B1",x"0C", -- 0x3B90
    x"4F",x"27",x"CC",x"8E",x"00",x"13",x"C6",x"04", -- 0x3B98
    x"D7",x"03",x"C6",x"01",x"96",x"50",x"91",x"5D", -- 0x3BA0
    x"26",x"13",x"96",x"51",x"91",x"5E",x"26",x"0D", -- 0x3BA8
    x"96",x"52",x"91",x"5F",x"26",x"07",x"96",x"53", -- 0x3BB0
    x"91",x"60",x"26",x"01",x"43",x"1F",x"A8",x"59", -- 0x3BB8
    x"24",x"0A",x"E7",x"80",x"0A",x"03",x"2B",x"34", -- 0x3BC0
    x"27",x"2E",x"C6",x"01",x"1F",x"8A",x"25",x"0E", -- 0x3BC8
    x"08",x"60",x"09",x"5F",x"09",x"5E",x"09",x"5D", -- 0x3BD0
    x"25",x"E3",x"2B",x"C8",x"20",x"DF",x"96",x"60", -- 0x3BD8
    x"90",x"53",x"97",x"60",x"96",x"5F",x"92",x"52", -- 0x3BE0
    x"97",x"5F",x"96",x"5E",x"92",x"51",x"97",x"5E", -- 0x3BE8
    x"96",x"5D",x"92",x"50",x"97",x"5D",x"20",x"D8", -- 0x3BF0
    x"C6",x"40",x"20",x"D0",x"56",x"56",x"56",x"D7", -- 0x3BF8
    x"63",x"8D",x"08",x"7E",x"BA",x"1C",x"C6",x"14", -- 0x3C00
    x"7E",x"AC",x"46",x"9E",x"13",x"9F",x"50",x"9E", -- 0x3C08
    x"15",x"9F",x"52",x"39",x"34",x"02",x"EC",x"01", -- 0x3C10
    x"97",x"54",x"8A",x"80",x"DD",x"50",x"0F",x"63", -- 0x3C18
    x"E6",x"84",x"AE",x"03",x"9F",x"52",x"D7",x"4F", -- 0x3C20
    x"35",x"82",x"8E",x"00",x"45",x"20",x"06",x"8E", -- 0x3C28
    x"00",x"40",x"8C",x"9E",x"3B",x"96",x"4F",x"A7", -- 0x3C30
    x"84",x"96",x"54",x"8A",x"7F",x"94",x"50",x"A7", -- 0x3C38
    x"01",x"96",x"51",x"A7",x"02",x"DE",x"52",x"EF", -- 0x3C40
    x"03",x"39",x"96",x"61",x"97",x"54",x"9E",x"5C", -- 0x3C48
    x"9F",x"4F",x"0F",x"63",x"96",x"5E",x"97",x"51", -- 0x3C50
    x"96",x"54",x"9E",x"5F",x"9F",x"52",x"39",x"DC", -- 0x3C58
    x"4F",x"DD",x"5C",x"9E",x"51",x"9F",x"5E",x"9E", -- 0x3C60
    x"53",x"9F",x"60",x"4D",x"39",x"D6",x"4F",x"27", -- 0x3C68
    x"08",x"D6",x"54",x"59",x"C6",x"FF",x"25",x"01", -- 0x3C70
    x"50",x"39",x"8D",x"F1",x"D7",x"50",x"0F",x"51", -- 0x3C78
    x"C6",x"88",x"96",x"50",x"80",x"80",x"D7",x"4F", -- 0x3C80
    x"DC",x"8A",x"DD",x"52",x"97",x"63",x"97",x"54", -- 0x3C88
    x"7E",x"BA",x"18",x"0F",x"54",x"39",x"E6",x"84", -- 0x3C90
    x"27",x"D3",x"E6",x"01",x"D8",x"54",x"2B",x"D1", -- 0x3C98
    x"D6",x"4F",x"E1",x"84",x"26",x"1D",x"E6",x"01", -- 0x3CA0
    x"CA",x"7F",x"D4",x"50",x"E1",x"01",x"26",x"13", -- 0x3CA8
    x"D6",x"51",x"E1",x"02",x"26",x"0D",x"D6",x"52", -- 0x3CB0
    x"E1",x"03",x"26",x"07",x"D6",x"53",x"E0",x"04", -- 0x3CB8
    x"26",x"01",x"39",x"56",x"D8",x"54",x"20",x"AB", -- 0x3CC0
    x"D6",x"4F",x"27",x"3D",x"C0",x"A0",x"96",x"54", -- 0x3CC8
    x"2A",x"05",x"03",x"5B",x"BD",x"BA",x"7B",x"8E", -- 0x3CD0
    x"00",x"4F",x"C1",x"F8",x"2E",x"06",x"BD",x"BA", -- 0x3CD8
    x"AE",x"0F",x"5B",x"39",x"0F",x"5B",x"96",x"54", -- 0x3CE0
    x"49",x"06",x"50",x"7E",x"BA",x"BA",x"D6",x"4F", -- 0x3CE8
    x"C1",x"A0",x"24",x"1D",x"8D",x"D2",x"D7",x"63", -- 0x3CF0
    x"96",x"54",x"D7",x"54",x"80",x"80",x"86",x"A0", -- 0x3CF8
    x"97",x"4F",x"96",x"53",x"97",x"01",x"7E",x"BA", -- 0x3D00
    x"18",x"D7",x"50",x"D7",x"51",x"D7",x"52",x"D7", -- 0x3D08
    x"53",x"39",x"9E",x"8A",x"9F",x"54",x"9F",x"4F", -- 0x3D10
    x"9F",x"51",x"9F",x"52",x"9F",x"47",x"9F",x"45", -- 0x3D18
    x"25",x"64",x"BD",x"01",x"97",x"81",x"2D",x"26", -- 0x3D20
    x"04",x"03",x"55",x"20",x"04",x"81",x"2B",x"26", -- 0x3D28
    x"04",x"9D",x"9F",x"25",x"51",x"81",x"2E",x"27", -- 0x3D30
    x"28",x"81",x"45",x"26",x"28",x"9D",x"9F",x"25", -- 0x3D38
    x"64",x"81",x"AC",x"27",x"0E",x"81",x"2D",x"27", -- 0x3D40
    x"0A",x"81",x"AB",x"27",x"08",x"81",x"2B",x"27", -- 0x3D48
    x"04",x"20",x"06",x"03",x"48",x"9D",x"9F",x"25", -- 0x3D50
    x"4C",x"0D",x"48",x"27",x"08",x"00",x"47",x"20", -- 0x3D58
    x"04",x"03",x"46",x"26",x"CC",x"96",x"47",x"90", -- 0x3D60
    x"45",x"97",x"47",x"27",x"12",x"2A",x"09",x"BD", -- 0x3D68
    x"BB",x"82",x"0C",x"47",x"26",x"F9",x"20",x"07", -- 0x3D70
    x"BD",x"BB",x"6A",x"0A",x"47",x"26",x"F9",x"96", -- 0x3D78
    x"55",x"2A",x"8E",x"7E",x"BE",x"E9",x"D6",x"45", -- 0x3D80
    x"D0",x"46",x"D7",x"45",x"34",x"02",x"BD",x"BB", -- 0x3D88
    x"6A",x"35",x"04",x"C0",x"30",x"8D",x"02",x"20", -- 0x3D90
    x"98",x"BD",x"BC",x"2F",x"BD",x"BC",x"7C",x"8E", -- 0x3D98
    x"00",x"40",x"7E",x"B9",x"C2",x"D6",x"47",x"58", -- 0x3DA0
    x"58",x"DB",x"47",x"58",x"80",x"30",x"34",x"04", -- 0x3DA8
    x"AB",x"E0",x"97",x"47",x"20",x"9F",x"9B",x"3E", -- 0x3DB0
    x"BC",x"1F",x"FD",x"9E",x"6E",x"6B",x"27",x"FD", -- 0x3DB8
    x"9E",x"6E",x"6B",x"28",x"00",x"8E",x"AB",x"E7", -- 0x3DC0
    x"8D",x"0C",x"DC",x"68",x"DD",x"50",x"C6",x"90", -- 0x3DC8
    x"43",x"BD",x"BC",x"86",x"8D",x"03",x"7E",x"B9", -- 0x3DD0
    x"9C",x"CE",x"03",x"DA",x"86",x"20",x"D6",x"54", -- 0x3DD8
    x"2A",x"02",x"86",x"2D",x"A7",x"C0",x"DF",x"64", -- 0x3DE0
    x"97",x"54",x"86",x"30",x"D6",x"4F",x"10",x"27", -- 0x3DE8
    x"00",x"C6",x"4F",x"C1",x"80",x"22",x"08",x"8E", -- 0x3DF0
    x"BD",x"C0",x"BD",x"BA",x"CA",x"86",x"F7",x"97", -- 0x3DF8
    x"45",x"8E",x"BD",x"BB",x"BD",x"BC",x"A0",x"2E", -- 0x3E00
    x"0F",x"8E",x"BD",x"B6",x"BD",x"BC",x"A0",x"2E", -- 0x3E08
    x"0E",x"BD",x"BB",x"6A",x"0A",x"45",x"20",x"F1", -- 0x3E10
    x"BD",x"BB",x"82",x"0C",x"45",x"20",x"E2",x"BD", -- 0x3E18
    x"B9",x"B4",x"BD",x"BC",x"C8",x"C6",x"01",x"96", -- 0x3E20
    x"45",x"8B",x"0A",x"2B",x"09",x"81",x"0B",x"24", -- 0x3E28
    x"05",x"4A",x"1F",x"89",x"86",x"02",x"4A",x"4A", -- 0x3E30
    x"97",x"47",x"D7",x"45",x"2E",x"0D",x"DE",x"64", -- 0x3E38
    x"86",x"2E",x"A7",x"C0",x"5D",x"27",x"04",x"86", -- 0x3E40
    x"30",x"A7",x"C0",x"8E",x"BE",x"C5",x"C6",x"80", -- 0x3E48
    x"96",x"53",x"AB",x"03",x"97",x"53",x"96",x"52", -- 0x3E50
    x"A9",x"02",x"97",x"52",x"96",x"51",x"A9",x"01", -- 0x3E58
    x"97",x"51",x"96",x"50",x"A9",x"84",x"97",x"50", -- 0x3E60
    x"5C",x"56",x"59",x"28",x"E3",x"24",x"03",x"C0", -- 0x3E68
    x"0B",x"50",x"CB",x"2F",x"30",x"04",x"1F",x"98", -- 0x3E70
    x"84",x"7F",x"A7",x"C0",x"0A",x"45",x"26",x"04", -- 0x3E78
    x"86",x"2E",x"A7",x"C0",x"53",x"C4",x"80",x"8C", -- 0x3E80
    x"BE",x"E9",x"26",x"C4",x"A6",x"C2",x"81",x"30", -- 0x3E88
    x"27",x"FA",x"81",x"2E",x"26",x"02",x"33",x"5F", -- 0x3E90
    x"86",x"2B",x"D6",x"47",x"27",x"1C",x"2A",x"03", -- 0x3E98
    x"86",x"2D",x"50",x"A7",x"42",x"86",x"45",x"A7", -- 0x3EA0
    x"41",x"86",x"2F",x"4C",x"C0",x"0A",x"24",x"FB", -- 0x3EA8
    x"CB",x"3A",x"ED",x"43",x"6F",x"45",x"20",x"04", -- 0x3EB0
    x"A7",x"C4",x"6F",x"41",x"8E",x"03",x"DA",x"39", -- 0x3EB8
    x"80",x"00",x"00",x"00",x"00",x"FA",x"0A",x"1F", -- 0x3EC0
    x"00",x"00",x"98",x"96",x"80",x"FF",x"F0",x"BD", -- 0x3EC8
    x"C0",x"00",x"01",x"86",x"A0",x"FF",x"FF",x"D8", -- 0x3ED0
    x"F0",x"00",x"00",x"03",x"E8",x"FF",x"FF",x"FF", -- 0x3ED8
    x"9C",x"00",x"00",x"00",x"0A",x"FF",x"FF",x"FF", -- 0x3EE0
    x"FF",x"96",x"4F",x"27",x"02",x"03",x"54",x"39", -- 0x3EE8
    x"9F",x"64",x"BD",x"BC",x"2F",x"8D",x"05",x"8D", -- 0x3EF0
    x"08",x"8E",x"00",x"40",x"7E",x"BA",x"CA",x"9F", -- 0x3EF8
    x"64",x"BD",x"BC",x"2A",x"9E",x"64",x"E6",x"80", -- 0x3F00
    x"D7",x"55",x"9F",x"64",x"8D",x"EE",x"9E",x"64", -- 0x3F08
    x"30",x"05",x"9F",x"64",x"BD",x"B9",x"C2",x"8E", -- 0x3F10
    x"00",x"45",x"0A",x"55",x"26",x"EE",x"39",x"BD", -- 0x3F18
    x"BC",x"6D",x"2B",x"21",x"27",x"15",x"8D",x"10", -- 0x3F20
    x"BD",x"BC",x"2F",x"8D",x"0E",x"8E",x"00",x"40", -- 0x3F28
    x"8D",x"CA",x"8E",x"BA",x"C5",x"BD",x"B9",x"C2", -- 0x3F30
    x"7E",x"BC",x"EE",x"BE",x"01",x"16",x"9F",x"50", -- 0x3F38
    x"BE",x"01",x"18",x"9F",x"52",x"BE",x"BF",x"74", -- 0x3F40
    x"9F",x"5D",x"BE",x"BF",x"76",x"9F",x"5F",x"BD", -- 0x3F48
    x"BA",x"D0",x"DC",x"AD",x"C3",x"65",x"8B",x"FD", -- 0x3F50
    x"01",x"18",x"DD",x"52",x"DC",x"AB",x"C9",x"B0", -- 0x3F58
    x"89",x"05",x"FD",x"01",x"16",x"DD",x"50",x"0F", -- 0x3F60
    x"54",x"86",x"80",x"97",x"4F",x"96",x"15",x"97", -- 0x3F68
    x"63",x"7E",x"BA",x"1C",x"40",x"E6",x"4D",x"AB", -- 0x3F70
    x"BD",x"BC",x"5F",x"8E",x"BF",x"BD",x"D6",x"61", -- 0x3F78
    x"BD",x"BB",x"89",x"BD",x"BC",x"5F",x"8D",x"B0", -- 0x3F80
    x"0F",x"62",x"96",x"5C",x"D6",x"4F",x"BD",x"B9", -- 0x3F88
    x"BC",x"8E",x"BF",x"C2",x"BD",x"B9",x"B9",x"96", -- 0x3F90
    x"54",x"34",x"02",x"2A",x"09",x"BD",x"B9",x"B4", -- 0x3F98
    x"96",x"54",x"2B",x"05",x"03",x"0A",x"BD",x"BE", -- 0x3FA0
    x"E9",x"8E",x"BF",x"C2",x"BD",x"B9",x"C2",x"35", -- 0x3FA8
    x"02",x"4D",x"2A",x"03",x"BD",x"BE",x"E9",x"8E", -- 0x3FB0
    x"BF",x"C7",x"7E",x"BE",x"F0",x"83",x"49",x"0F", -- 0x3FB8
    x"DA",x"A2",x"7F",x"00",x"00",x"00",x"00",x"05", -- 0x3FC0
    x"84",x"E6",x"1A",x"2D",x"1B",x"86",x"28",x"07", -- 0x3FC8
    x"FB",x"F8",x"87",x"99",x"68",x"89",x"01",x"87", -- 0x3FD0
    x"23",x"35",x"DF",x"E1",x"86",x"A5",x"5D",x"E7", -- 0x3FD8
    x"28",x"83",x"49",x"0F",x"DA",x"A2",x"A1",x"54", -- 0x3FE0
    x"46",x"8F",x"13",x"8F",x"52",x"43",x"89",x"CD", -- 0x3FE8
    x"A6",x"81",x"FE",x"EE",x"FE",x"F1",x"FE",x"F4", -- 0x3FF0
    x"FE",x"F7",x"FE",x"FA",x"FE",x"FD",x"8C",x"1B", -- 0x3FF8
    x"1A",x"50",x"10",x"CE",x"5E",x"FF",x"86",x"12", -- 0x4000
    x"C6",x"10",x"8E",x"FF",x"B0",x"A7",x"80",x"5A", -- 0x4008
    x"26",x"FB",x"8E",x"FF",x"A0",x"31",x"8D",x"02", -- 0x4010
    x"2D",x"C6",x"10",x"A6",x"A0",x"A7",x"80",x"5A", -- 0x4018
    x"26",x"F9",x"86",x"CE",x"B7",x"FF",x"90",x"30", -- 0x4020
    x"8D",x"00",x"14",x"10",x"8E",x"40",x"00",x"EC", -- 0x4028
    x"81",x"EE",x"81",x"ED",x"A1",x"EF",x"A1",x"8C", -- 0x4030
    x"C3",x"6C",x"25",x"F3",x"7E",x"40",x"00",x"32", -- 0x4038
    x"7F",x"12",x"12",x"12",x"12",x"12",x"86",x"FF", -- 0x4040
    x"B7",x"FF",x"94",x"B7",x"FF",x"95",x"30",x"8D", -- 0x4048
    x"01",x"DC",x"10",x"8E",x"FF",x"98",x"A6",x"80", -- 0x4050
    x"A7",x"A0",x"10",x"8C",x"FF",x"A0",x"26",x"F6", -- 0x4058
    x"8E",x"FF",x"20",x"CC",x"FF",x"34",x"6F",x"01", -- 0x4060
    x"6F",x"03",x"4A",x"A7",x"84",x"86",x"F8",x"A7", -- 0x4068
    x"02",x"E7",x"01",x"E7",x"03",x"6F",x"02",x"86", -- 0x4070
    x"02",x"A7",x"84",x"86",x"FF",x"8E",x"FF",x"00", -- 0x4078
    x"6F",x"01",x"6F",x"03",x"6F",x"84",x"A7",x"02", -- 0x4080
    x"E7",x"01",x"E7",x"03",x"C6",x"0C",x"CE",x"FF", -- 0x4088
    x"C0",x"A7",x"C1",x"5A",x"26",x"FB",x"B7",x"FF", -- 0x4090
    x"C9",x"1F",x"9B",x"6F",x"02",x"A7",x"5D",x"8E", -- 0x4098
    x"FF",x"00",x"C6",x"DF",x"E7",x"02",x"A6",x"84", -- 0x40A0
    x"43",x"84",x"40",x"A7",x"E4",x"10",x"8E",x"00", -- 0x40A8
    x"02",x"57",x"E7",x"02",x"A6",x"84",x"43",x"84", -- 0x40B0
    x"40",x"27",x"07",x"31",x"3F",x"26",x"F2",x"16", -- 0x40B8
    x"01",x"2E",x"86",x"CA",x"B7",x"FF",x"90",x"B6", -- 0x40C0
    x"FE",x"ED",x"81",x"55",x"26",x"28",x"96",x"71", -- 0x40C8
    x"81",x"55",x"26",x"0A",x"9E",x"72",x"A6",x"84", -- 0x40D0
    x"81",x"12",x"10",x"27",x"00",x"AE",x"7F",x"FF", -- 0x40D8
    x"A0",x"96",x"71",x"81",x"55",x"26",x"0A",x"9E", -- 0x40E0
    x"72",x"A6",x"84",x"81",x"12",x"10",x"27",x"00", -- 0x40E8
    x"9B",x"86",x"38",x"B7",x"FF",x"A0",x"8E",x"C0", -- 0x40F0
    x"00",x"10",x"8E",x"80",x"00",x"17",x"00",x"AA", -- 0x40F8
    x"31",x"8D",x"01",x"52",x"A6",x"A0",x"34",x"02", -- 0x4100
    x"AE",x"A1",x"E6",x"A0",x"A6",x"A0",x"A7",x"80", -- 0x4108
    x"5A",x"26",x"F9",x"35",x"02",x"4A",x"26",x"EE", -- 0x4110
    x"7F",x"FF",x"DE",x"86",x"C8",x"B7",x"FF",x"90", -- 0x4118
    x"FC",x"C0",x"00",x"81",x"44",x"26",x"10",x"C1", -- 0x4120
    x"4B",x"26",x"0C",x"8E",x"E0",x"00",x"10",x"8E", -- 0x4128
    x"C0",x"00",x"8D",x"76",x"17",x"01",x"EB",x"7F", -- 0x4130
    x"FF",x"DE",x"86",x"CA",x"B7",x"FF",x"90",x"8E", -- 0x4138
    x"FE",x"00",x"10",x"8E",x"E0",x"00",x"8D",x"62", -- 0x4140
    x"17",x"00",x"93",x"31",x"8D",x"02",x"0A",x"8E", -- 0x4148
    x"FE",x"ED",x"C6",x"13",x"17",x"00",x"7F",x"7F", -- 0x4150
    x"FF",x"DF",x"6D",x"E4",x"27",x"22",x"8E",x"E0", -- 0x4158
    x"32",x"C6",x"03",x"30",x"01",x"A6",x"84",x"8A", -- 0x4160
    x"20",x"A7",x"84",x"30",x"09",x"5A",x"26",x"F5", -- 0x4168
    x"C6",x"02",x"8E",x"E0",x"70",x"A6",x"84",x"8A", -- 0x4170
    x"20",x"A7",x"84",x"30",x"09",x"5A",x"26",x"F5", -- 0x4178
    x"8E",x"04",x"00",x"86",x"60",x"A7",x"80",x"8C", -- 0x4180
    x"06",x"00",x"25",x"F9",x"86",x"CE",x"B7",x"FF", -- 0x4188
    x"90",x"6D",x"E4",x"27",x"05",x"86",x"20",x"B7", -- 0x4190
    x"FF",x"98",x"8E",x"FF",x"B0",x"31",x"8D",x"00", -- 0x4198
    x"95",x"C6",x"10",x"8D",x"31",x"32",x"61",x"7E", -- 0x41A0
    x"A0",x"27",x"BF",x"5F",x"02",x"10",x"FF",x"5F", -- 0x41A8
    x"00",x"7F",x"FF",x"DE",x"EC",x"A4",x"AE",x"22", -- 0x41B0
    x"EE",x"24",x"10",x"EE",x"26",x"7F",x"FF",x"DF", -- 0x41B8
    x"ED",x"A4",x"AF",x"22",x"EF",x"24",x"10",x"EF", -- 0x41C0
    x"26",x"31",x"28",x"10",x"BC",x"5F",x"02",x"25", -- 0x41C8
    x"E0",x"10",x"FE",x"5F",x"00",x"39",x"A6",x"A0", -- 0x41D0
    x"A7",x"80",x"5A",x"26",x"F9",x"39",x"8E",x"F7", -- 0x41D8
    x"1B",x"31",x"8D",x"01",x"28",x"C6",x"15",x"A6", -- 0x41E0
    x"A0",x"43",x"A7",x"80",x"5A",x"26",x"F8",x"39", -- 0x41E8
    x"4F",x"B7",x"FE",x"ED",x"97",x"71",x"B7",x"FF", -- 0x41F0
    x"DE",x"C6",x"09",x"F7",x"FF",x"BA",x"C6",x"3F", -- 0x41F8
    x"F7",x"FF",x"BB",x"8E",x"C4",x"05",x"10",x"8E", -- 0x4200
    x"0E",x"00",x"EC",x"81",x"EE",x"81",x"ED",x"A1", -- 0x4208
    x"EF",x"A1",x"8C",x"DC",x"05",x"25",x"F3",x"86", -- 0x4210
    x"F9",x"B7",x"FF",x"22",x"4F",x"8E",x"FF",x"C0", -- 0x4218
    x"A7",x"84",x"A7",x"03",x"A7",x"05",x"A7",x"07", -- 0x4220
    x"A7",x"09",x"A7",x"0B",x"20",x"FE",x"00",x"00", -- 0x4228
    x"00",x"00",x"0F",x"E0",x"00",x"00",x"12",x"24", -- 0x4230
    x"0B",x"07",x"3F",x"1F",x"09",x"26",x"00",x"12", -- 0x4238
    x"00",x"3F",x"00",x"12",x"00",x"26",x"38",x"39", -- 0x4240
    x"34",x"3B",x"3C",x"3D",x"3E",x"3F",x"38",x"30", -- 0x4248
    x"31",x"32",x"33",x"3D",x"35",x"3F",x"1B",x"80", -- 0x4250
    x"C0",x"01",x"12",x"B8",x"D4",x"03",x"7E",x"E1", -- 0x4258
    x"38",x"B7",x"F3",x"03",x"7E",x"E1",x"72",x"81", -- 0x4260
    x"50",x"04",x"7E",x"E1",x"92",x"12",x"81",x"6C", -- 0x4268
    x"04",x"7E",x"E1",x"A6",x"12",x"88",x"34",x"12", -- 0x4270
    x"7E",x"E3",x"F8",x"0F",x"51",x"0F",x"52",x"0F", -- 0x4278
    x"53",x"20",x"B0",x"0F",x"50",x"20",x"CF",x"7E", -- 0x4280
    x"E4",x"0C",x"87",x"EB",x"07",x"20",x"4A",x"12", -- 0x4288
    x"39",x"8E",x"00",x"51",x"88",x"0C",x"02",x"20", -- 0x4290
    x"35",x"88",x"26",x"02",x"25",x"17",x"87",x"E7", -- 0x4298
    x"02",x"26",x"05",x"88",x"6A",x"02",x"26",x"82", -- 0x42A0
    x"80",x"B2",x"03",x"7E",x"E2",x"88",x"81",x"3A", -- 0x42A8
    x"01",x"00",x"97",x"03",x"03",x"7E",x"E3",x"89", -- 0x42B0
    x"AD",x"F0",x"04",x"7E",x"E4",x"29",x"12",x"A3", -- 0x42B8
    x"C2",x"04",x"7E",x"E4",x"13",x"12",x"B0",x"3D", -- 0x42C0
    x"02",x"E5",x"32",x"AF",x"42",x"03",x"7E",x"E3", -- 0x42C8
    x"B4",x"AD",x"3F",x"04",x"7E",x"E4",x"D0",x"12", -- 0x42D0
    x"AC",x"46",x"03",x"7E",x"E4",x"70",x"AC",x"73", -- 0x42D8
    x"03",x"7E",x"E5",x"02",x"A3",x"0A",x"03",x"7E", -- 0x42E0
    x"8C",x"37",x"A9",x"10",x"03",x"7E",x"8C",x"46", -- 0x42E8
    x"A1",x"B1",x"08",x"7E",x"A0",x"CE",x"12",x"12", -- 0x42F0
    x"12",x"12",x"12",x"B9",x"02",x"03",x"7E",x"F8", -- 0x42F8
    x"C3",x"B9",x"5C",x"03",x"7E",x"F8",x"A3",x"A3", -- 0x4300
    x"8D",x"03",x"7E",x"F7",x"57",x"AB",x"D1",x"B7", -- 0x4308
    x"9E",x"8D",x"8D",x"96",x"8C",x"DF",x"D9",x"DF", -- 0x4310
    x"AB",x"D1",x"BA",x"9E",x"8D",x"93",x"9A",x"8C", -- 0x4318
    x"F2",x"FF",x"B6",x"C0",x"04",x"81",x"D6",x"26", -- 0x4320
    x"0B",x"8E",x"C0",x"C6",x"31",x"8D",x"00",x"25", -- 0x4328
    x"E6",x"A0",x"20",x"15",x"8E",x"C8",x"B4",x"86", -- 0x4330
    x"12",x"C6",x"0B",x"A7",x"80",x"5A",x"26",x"FB", -- 0x4338
    x"8E",x"C0",x"D9",x"31",x"8D",x"00",x"0A",x"E6", -- 0x4340
    x"A0",x"A6",x"A0",x"A7",x"80",x"5A",x"26",x"F9", -- 0x4348
    x"39",x"03",x"7E",x"E2",x"9D",x"03",x"7E",x"E2", -- 0x4350
    x"97",x"55",x"16",x"02",x"0F",x"16",x"02",x"0F", -- 0x4358
    x"16",x"02",x"18",x"16",x"02",x"12",x"16",x"02", -- 0x4360
    x"09",x"16",x"02",x"09",x"FF",x"FF",x"FF",x"FF", -- 0x4368
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x4370
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4378
    x"00",x"55",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x4380
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4388
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x4390
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4398
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x43A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x43A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x43B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x43B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x43C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x43C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x43D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x43D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x43E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x43E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x43F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x43F8
    x"00",x"18",x"00",x"0E",x"00",x"FF",x"FF",x"FF", -- 0x4400
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4408
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4410
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4418
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4420
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4428
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4430
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4438
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4440
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4448
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4450
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4458
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4460
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4468
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4470
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4478
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4480
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4488
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4490
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4498
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x44A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x44A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x44B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x44B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x44C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x44C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x44D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x44D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"00", -- 0x44E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x44E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x44F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x44F8
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x4500
    x"FB",x"EE",x"EF",x"FB",x"FF",x"BB",x"FF",x"FF", -- 0x4508
    x"FF",x"FB",x"FF",x"FF",x"BB",x"BB",x"BB",x"BF", -- 0x4510
    x"BB",x"BB",x"FF",x"BF",x"FF",x"FE",x"EF",x"FF", -- 0x4518
    x"FF",x"FF",x"EF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4520
    x"FF",x"BB",x"BB",x"BF",x"FF",x"FF",x"FF",x"FF", -- 0x4528
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4530
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"BF", -- 0x4538
    x"BB",x"FF",x"BB",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4540
    x"EE",x"EE",x"EE",x"EE",x"EF",x"FF",x"FE",x"FF", -- 0x4548
    x"FE",x"EE",x"EE",x"FE",x"EE",x"EE",x"EE",x"EF", -- 0x4550
    x"EE",x"EE",x"EE",x"EE",x"EE",x"FE",x"EE",x"EE", -- 0x4558
    x"EE",x"EE",x"EE",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x4560
    x"FF",x"BB",x"BB",x"BB",x"BB",x"BF",x"FF",x"FF", -- 0x4568
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4570
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"BB",x"BB", -- 0x4578
    x"BB",x"BB",x"BB",x"7F",x"FF",x"FF",x"F6",x"AA", -- 0x4580
    x"AE",x"AA",x"AE",x"AA",x"EA",x"BB",x"BB",x"FB", -- 0x4588
    x"FF",x"BB",x"FF",x"BF",x"BF",x"FF",x"FB",x"BF", -- 0x4590
    x"BB",x"BB",x"BB",x"BB",x"BB",x"BA",x"EA",x"AA", -- 0x4598
    x"EE",x"AE",x"EE",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x45A0
    x"BF",x"BB",x"BB",x"BB",x"BB",x"BF",x"FF",x"FF", -- 0x45A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x45B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"BB",x"BB", -- 0x45B8
    x"BB",x"BB",x"BB",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x45C0
    x"EE",x"EE",x"EE",x"EE",x"EE",x"EE",x"EE",x"EF", -- 0x45C8
    x"FE",x"EF",x"FF",x"FF",x"FF",x"FF",x"FE",x"EF", -- 0x45D0
    x"EE",x"EE",x"EE",x"EE",x"EE",x"EE",x"EE",x"EE", -- 0x45D8
    x"EE",x"EE",x"EF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x45E0
    x"BB",x"BB",x"BB",x"BB",x"BB",x"BF",x"FF",x"FF", -- 0x45E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x45F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"BB", -- 0x45F8
    x"BB",x"BB",x"BB",x"7F",x"FF",x"FF",x"F6",x"AA", -- 0x4600
    x"EE",x"AA",x"AA",x"AA",x"EA",x"AB",x"BB",x"BB", -- 0x4608
    x"FF",x"BB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4610
    x"FB",x"BF",x"FF",x"FF",x"BB",x"BB",x"EA",x"AE", -- 0x4618
    x"AA",x"AA",x"AF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4620
    x"BB",x"BF",x"FF",x"FB",x"BB",x"BF",x"FF",x"FF", -- 0x4628
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4630
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"BB", -- 0x4638
    x"BB",x"BB",x"BB",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4640
    x"EE",x"EE",x"EF",x"EF",x"EE",x"EE",x"EF",x"FF", -- 0x4648
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4650
    x"FF",x"FF",x"FF",x"FF",x"EE",x"EE",x"FF",x"EF", -- 0x4658
    x"EE",x"EE",x"EF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4660
    x"BB",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4668
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4670
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4678
    x"BB",x"BB",x"BB",x"7F",x"FF",x"FF",x"F7",x"EA", -- 0x4680
    x"AA",x"BB",x"BB",x"BB",x"BB",x"BB",x"FB",x"BB", -- 0x4688
    x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4690
    x"FF",x"FB",x"FF",x"FB",x"FB",x"BB",x"BB",x"BA", -- 0x4698
    x"AA",x"AA",x"EF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x46A0
    x"BB",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x46A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x46B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB", -- 0x46B8
    x"BB",x"BB",x"BB",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x46C0
    x"EE",x"EE",x"FE",x"EE",x"EE",x"EE",x"EE",x"FF", -- 0x46C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x46D0
    x"FF",x"FF",x"FF",x"FE",x"EE",x"EF",x"FE",x"EE", -- 0x46D8
    x"EE",x"EE",x"EF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x46E0
    x"BB",x"FB",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x46E8
    x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x46F0
    x"00",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB", -- 0x46F8
    x"BB",x"BB",x"BB",x"7F",x"FF",x"FF",x"F6",x"EA", -- 0x4700
    x"AB",x"AA",x"AB",x"BB",x"BB",x"BF",x"BF",x"FF", -- 0x4708
    x"FF",x"FF",x"80",x"00",x"7F",x"FF",x"FF",x"C0", -- 0x4710
    x"00",x"3F",x"FF",x"FF",x"BB",x"BB",x"BF",x"AA", -- 0x4718
    x"AA",x"AA",x"EF",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x4720
    x"BB",x"BB",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4728
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4730
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BB", -- 0x4738
    x"BB",x"BB",x"BF",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4740
    x"EE",x"EE",x"EF",x"EE",x"FF",x"FF",x"FF",x"EE", -- 0x4748
    x"FF",x"FF",x"80",x"00",x"3F",x"FF",x"FF",x"80", -- 0x4750
    x"00",x"3F",x"FF",x"FF",x"EE",x"FE",x"EE",x"EE", -- 0x4758
    x"EE",x"EE",x"EF",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x4760
    x"BB",x"BB",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4768
    x"FF",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x4770
    x"00",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",x"BB", -- 0x4778
    x"BB",x"BB",x"BF",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4780
    x"AB",x"AE",x"EB",x"BB",x"BF",x"FB",x"FF",x"FF", -- 0x4788
    x"FF",x"FF",x"80",x"00",x"1F",x"FF",x"FF",x"00", -- 0x4790
    x"00",x"3F",x"FF",x"FF",x"FF",x"BB",x"BB",x"AA", -- 0x4798
    x"AA",x"BE",x"AB",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x47A0
    x"BF",x"BB",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x47A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x47B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FB", -- 0x47B8
    x"BB",x"BB",x"BF",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x47C0
    x"EE",x"EE",x"EE",x"EE",x"EF",x"FE",x"EF",x"FF", -- 0x47C8
    x"FF",x"FF",x"80",x"00",x"0F",x"FF",x"FE",x"00", -- 0x47D0
    x"00",x"3F",x"FF",x"FF",x"EF",x"EF",x"EE",x"EE", -- 0x47D8
    x"EE",x"EE",x"EF",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x47E0
    x"BF",x"FB",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x47E8
    x"FF",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x47F0
    x"00",x"03",x"FF",x"FF",x"FF",x"FF",x"FB",x"BF", -- 0x47F8
    x"FF",x"BB",x"BF",x"7F",x"FF",x"FF",x"F6",x"EA", -- 0x4800
    x"AB",x"BA",x"AB",x"BB",x"FB",x"FF",x"BF",x"FF", -- 0x4808
    x"FF",x"FF",x"80",x"00",x"07",x"FF",x"FC",x"00", -- 0x4810
    x"00",x"3F",x"FF",x"FF",x"FF",x"FB",x"AA",x"FF", -- 0x4818
    x"FE",x"EA",x"AB",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x4820
    x"BF",x"FB",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4828
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4830
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"BF", -- 0x4838
    x"FF",x"BB",x"BF",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4840
    x"EE",x"FF",x"FE",x"EE",x"EE",x"FF",x"FF",x"FF", -- 0x4848
    x"FF",x"FF",x"80",x"00",x"03",x"FF",x"F8",x"00", -- 0x4850
    x"00",x"3F",x"FF",x"FF",x"FE",x"EE",x"EE",x"FF", -- 0x4858
    x"FE",x"EE",x"EF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4860
    x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4868
    x"FF",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x4870
    x"00",x"03",x"FF",x"FF",x"FF",x"FF",x"BB",x"BF", -- 0x4878
    x"FF",x"BB",x"FF",x"7F",x"FF",x"FF",x"F7",x"AA", -- 0x4880
    x"FB",x"BB",x"BB",x"BF",x"FF",x"FF",x"FF",x"FF", -- 0x4888
    x"FF",x"FF",x"80",x"00",x"01",x"FF",x"F0",x"00", -- 0x4890
    x"00",x"3F",x"FF",x"FF",x"BB",x"BB",x"AE",x"BB", -- 0x4898
    x"BE",x"AF",x"BB",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x48A0
    x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x48A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x48B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"FF", -- 0x48B8
    x"FF",x"BB",x"FF",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x48C0
    x"EE",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF", -- 0x48C8
    x"FF",x"FF",x"80",x"08",x"00",x"FF",x"E0",x"02", -- 0x48D0
    x"00",x"3F",x"FF",x"FF",x"FE",x"EF",x"EE",x"FF", -- 0x48D8
    x"EE",x"EF",x"EF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x48E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x48E8
    x"FF",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x48F0
    x"00",x"03",x"FF",x"FF",x"FF",x"FF",x"FB",x"FF", -- 0x48F8
    x"FF",x"BB",x"FF",x"7F",x"FF",x"FF",x"F7",x"AA", -- 0x4900
    x"BB",x"BB",x"FB",x"BB",x"FF",x"BF",x"FF",x"FF", -- 0x4908
    x"FF",x"FF",x"80",x"0C",x"00",x"7F",x"C0",x"06", -- 0x4910
    x"00",x"3F",x"FF",x"FF",x"FF",x"BB",x"FF",x"FF", -- 0x4918
    x"BF",x"EB",x"BB",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4920
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4928
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4930
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4938
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4940
    x"EF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4948
    x"FF",x"FF",x"80",x"0E",x"00",x"3F",x"80",x"0E", -- 0x4950
    x"00",x"3F",x"FF",x"FF",x"FE",x"FF",x"FF",x"FE", -- 0x4958
    x"EE",x"EE",x"FF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4960
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4968
    x"FF",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x4970
    x"00",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4978
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F3",x"EA", -- 0x4980
    x"BB",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4988
    x"FF",x"FF",x"80",x"0F",x"00",x"1F",x"00",x"1E", -- 0x4990
    x"00",x"3F",x"FF",x"FF",x"FF",x"BF",x"FF",x"FF", -- 0x4998
    x"FF",x"FF",x"BF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x49A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x49A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x49B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x49B8
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"EE", -- 0x49C0
    x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x49C8
    x"FF",x"FF",x"80",x"0F",x"80",x"0E",x"00",x"3E", -- 0x49D0
    x"00",x"3F",x"FF",x"FF",x"EE",x"FF",x"FF",x"FF", -- 0x49D8
    x"FE",x"EF",x"EF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x49E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x49E8
    x"FF",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x49F0
    x"00",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x49F8
    x"FF",x"FF",x"BF",x"7F",x"FF",x"FF",x"F6",x"EA", -- 0x4A00
    x"BB",x"BB",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4A08
    x"FF",x"FF",x"80",x"0F",x"C0",x"00",x"00",x"7E", -- 0x4A10
    x"00",x"3F",x"FF",x"FF",x"BF",x"FF",x"FF",x"FF", -- 0x4A18
    x"FF",x"BA",x"EF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4A20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4A28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"1F",x"FF", -- 0x4A30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4A38
    x"FF",x"FF",x"BB",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4A40
    x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4A48
    x"FF",x"FF",x"80",x"0F",x"E0",x"00",x"00",x"FE", -- 0x4A50
    x"00",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4A58
    x"FE",x"FE",x"EF",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4A60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4A68
    x"FF",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x4A70
    x"00",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4A78
    x"FF",x"FF",x"BB",x"7F",x"FF",x"FF",x"F6",x"EB", -- 0x4A80
    x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4A88
    x"FF",x"FF",x"80",x"0F",x"C0",x"00",x"00",x"3E", -- 0x4A90
    x"00",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4A98
    x"FF",x"FE",x"EB",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4AA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4AA8
    x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"1F", -- 0x4AB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4AB8
    x"FF",x"FF",x"BA",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4AC0
    x"EF",x"FF",x"FF",x"FF",x"C0",x"1F",x"FF",x"FF", -- 0x4AC8
    x"FF",x"FF",x"80",x"0C",x"00",x"00",x"00",x"1E", -- 0x4AD0
    x"00",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4AD8
    x"FF",x"EE",x"EB",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4AE0
    x"FF",x"FF",x"FF",x"FC",x"00",x"0F",x"FF",x"FF", -- 0x4AE8
    x"FF",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x4AF0
    x"00",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x4AF8
    x"FF",x"FE",x"AA",x"7F",x"FF",x"FF",x"F6",x"AB", -- 0x4B00
    x"BB",x"FF",x"FF",x"00",x"00",x"03",x"FF",x"FF", -- 0x4B08
    x"FF",x"FF",x"80",x"0C",x"00",x"00",x"00",x"06", -- 0x4B10
    x"00",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"79", -- 0x4B18
    x"9F",x"FB",x"AB",x"7F",x"FF",x"FF",x"F7",x"BB", -- 0x4B20
    x"FF",x"FF",x"F8",x"00",x"00",x"01",x"FF",x"FF", -- 0x4B28
    x"FF",x"FF",x"FF",x"F0",x"00",x"00",x"38",x"03", -- 0x4B30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"00", -- 0x4B38
    x"03",x"FE",x"EE",x"7F",x"FF",x"FF",x"F6",x"EF", -- 0x4B40
    x"FF",x"FF",x"E0",x"00",x"00",x"00",x"4F",x"FF", -- 0x4B48
    x"FF",x"FF",x"80",x"00",x"00",x"01",x"7C",x"00", -- 0x4B50
    x"00",x"3F",x"FF",x"FF",x"FF",x"FF",x"80",x"00", -- 0x4B58
    x"00",x"FA",x"BB",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x4B60
    x"FF",x"FF",x"C0",x"00",x"00",x"00",x"01",x"FF", -- 0x4B68
    x"FF",x"F0",x"00",x"00",x"00",x"03",x"FE",x"00", -- 0x4B70
    x"00",x"03",x"FF",x"FF",x"FF",x"FF",x"00",x"00", -- 0x4B78
    x"00",x"7E",x"EE",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x4B80
    x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF", -- 0x4B88
    x"FF",x"FF",x"80",x"00",x"00",x"0F",x"FF",x"00", -- 0x4B90
    x"00",x"3F",x"FF",x"FF",x"FF",x"FC",x"00",x"00", -- 0x4B98
    x"00",x"3B",x"BB",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x4BA0
    x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",x"7F", -- 0x4BA8
    x"FF",x"FF",x"FF",x"00",x"00",x"2F",x"FF",x"00", -- 0x4BB0
    x"7F",x"FF",x"FF",x"FF",x"FF",x"F0",x"00",x"00", -- 0x4BB8
    x"00",x"0E",x"EE",x"7F",x"FF",x"FF",x"F6",x"FF", -- 0x4BC0
    x"FF",x"FC",x"00",x"00",x"00",x"00",x"00",x"3F", -- 0x4BC8
    x"FF",x"FF",x"80",x"00",x"01",x"FF",x"FF",x"80", -- 0x4BD0
    x"00",x"3F",x"FF",x"FF",x"FF",x"E0",x"00",x"00", -- 0x4BD8
    x"00",x"07",x"BB",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x4BE0
    x"FF",x"F8",x"00",x"00",x"00",x"00",x"00",x"3F", -- 0x4BE8
    x"FF",x"F0",x"00",x"00",x"03",x"FF",x"FF",x"40", -- 0x4BF0
    x"00",x"03",x"FF",x"FF",x"FF",x"C0",x"00",x"00", -- 0x4BF8
    x"00",x"03",x"EE",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x4C00
    x"FF",x"F0",x"00",x"00",x"00",x"01",x"00",x"1F", -- 0x4C08
    x"FF",x"FF",x"80",x"01",x"07",x"FF",x"FF",x"A0", -- 0x4C10
    x"00",x"3F",x"FF",x"FF",x"FF",x"80",x"00",x"00", -- 0x4C18
    x"00",x"01",x"BB",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x4C20
    x"FF",x"E0",x"00",x"00",x"00",x"01",x"80",x"1F", -- 0x4C28
    x"FF",x"FF",x"FE",x"0E",x"2F",x"FF",x"FF",x"C0", -- 0x4C30
    x"1F",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00", -- 0x4C38
    x"00",x"00",x"EE",x"7F",x"FF",x"FF",x"F6",x"FF", -- 0x4C40
    x"FF",x"E0",x"00",x"00",x"00",x"65",x"E0",x"0F", -- 0x4C48
    x"FF",x"FF",x"80",x"0C",x"1F",x"FF",x"FF",x"E0", -- 0x4C50
    x"00",x"3F",x"FF",x"FF",x"FF",x"00",x"00",x"00", -- 0x4C58
    x"00",x"00",x"3B",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x4C60
    x"FF",x"C0",x"00",x"00",x"0B",x"FF",x"F0",x"0F", -- 0x4C68
    x"FF",x"FC",x"00",x"18",x"0F",x"F8",x"00",x"60", -- 0x4C70
    x"00",x"07",x"FF",x"FF",x"FE",x"00",x"00",x"00", -- 0x4C78
    x"00",x"00",x"0E",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x4C80
    x"FF",x"C0",x"00",x"01",x"FF",x"FF",x"F8",x"0F", -- 0x4C88
    x"FF",x"FF",x"80",x"00",x"01",x"F8",x"00",x"20", -- 0x4C90
    x"00",x"3F",x"FF",x"FF",x"FE",x"00",x"00",x"00", -- 0x4C98
    x"00",x"00",x"1B",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x4CA0
    x"FF",x"80",x"00",x"03",x"FF",x"FF",x"FC",x"0F", -- 0x4CA8
    x"FF",x"FF",x"FC",x"03",x"03",x"FF",x"7F",x"F0", -- 0x4CB0
    x"03",x"FF",x"FF",x"FF",x"FC",x"00",x"00",x"00", -- 0x4CB8
    x"00",x"00",x"0E",x"7F",x"FF",x"FF",x"F7",x"FE", -- 0x4CC0
    x"FF",x"80",x"01",x"5D",x"FF",x"FF",x"FC",x"0F", -- 0x4CC8
    x"FF",x"FF",x"C0",x"07",x"F1",x"FC",x"07",x"FC", -- 0x4CD0
    x"00",x"3F",x"FF",x"FF",x"FC",x"00",x"00",x"00", -- 0x4CD8
    x"00",x"00",x"03",x"7F",x"FF",x"FF",x"F7",x"BF", -- 0x4CE0
    x"FF",x"00",x"02",x"EF",x"FF",x"FF",x"FC",x"0F", -- 0x4CE8
    x"FF",x"FF",x"00",x"0E",x"00",x"7C",x"00",x"F4", -- 0x4CF0
    x"00",x"0C",x"7F",x"FF",x"F8",x"00",x"00",x"00", -- 0x4CF8
    x"00",x"00",x"0E",x"7F",x"FF",x"FF",x"F2",x"AB", -- 0x4D00
    x"FF",x"00",x"05",x"FF",x"FF",x"FF",x"FE",x"0F", -- 0x4D08
    x"FF",x"FF",x"F8",x"1C",x"00",x"FC",x"01",x"F8", -- 0x4D10
    x"01",x"FB",x"BF",x"FF",x"F8",x"00",x"00",x"0F", -- 0x4D18
    x"E1",x"80",x"0B",x"7F",x"FF",x"FF",x"F7",x"BF", -- 0x4D20
    x"FF",x"00",x"03",x"FF",x"FF",x"FF",x"FE",x"0F", -- 0x4D28
    x"FF",x"FF",x"F8",x"1F",x"C0",x"FE",x"3F",x"FC", -- 0x4D30
    x"01",x"F6",x"DF",x"FF",x"F8",x"00",x"3F",x"FF", -- 0x4D38
    x"FF",x"80",x"0E",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4D40
    x"EE",x"00",x"07",x"FF",x"FF",x"FF",x"FE",x"0F", -- 0x4D48
    x"FE",x"FF",x"FC",x"1F",x"F1",x"FF",x"9F",x"F8", -- 0x4D50
    x"37",x"F5",x"DF",x"FF",x"F8",x"00",x"FF",x"FF", -- 0x4D58
    x"FF",x"80",x"0B",x"7F",x"FF",x"FF",x"F7",x"BF", -- 0x4D60
    x"FF",x"00",x"07",x"FF",x"FF",x"FF",x"FF",x"07", -- 0x4D68
    x"FF",x"FF",x"F8",x"0F",x"EF",x"7F",x"FF",x"FC", -- 0x4D70
    x"03",x"F6",x"DF",x"FF",x"F8",x"7F",x"FF",x"FF", -- 0x4D78
    x"FF",x"80",x"06",x"7F",x"FF",x"FF",x"F6",x"FF", -- 0x4D80
    x"BF",x"00",x"03",x"FF",x"FF",x"FF",x"FF",x"07", -- 0x4D88
    x"FB",x"BB",x"FD",x"DF",x"FF",x"EF",x"FF",x"F9", -- 0x4D90
    x"7F",x"FB",x"BF",x"FF",x"FC",x"7F",x"FF",x"FF", -- 0x4D98
    x"FF",x"C0",x"0B",x"7F",x"FF",x"FF",x"F7",x"BF", -- 0x4DA0
    x"FE",x"00",x"03",x"FF",x"FF",x"FF",x"F8",x"07", -- 0x4DA8
    x"FF",x"FF",x"FF",x"9F",x"FF",x"FF",x"FF",x"FF", -- 0x4DB0
    x"BF",x"FC",x"7F",x"FF",x"FC",x"75",x"0F",x"FF", -- 0x4DB8
    x"CF",x"C0",x"0E",x"7F",x"FF",x"FF",x"F6",x"FF", -- 0x4DC0
    x"FE",x"00",x"07",x"F5",x"47",x"FF",x"E0",x"07", -- 0x4DC8
    x"FF",x"EF",x"FF",x"CF",x"FD",x"FF",x"FF",x"FF", -- 0x4DD0
    x"3F",x"FF",x"FF",x"FF",x"FC",x"00",x"00",x"E0", -- 0x4DD8
    x"07",x"C0",x"0F",x"7F",x"FF",x"FF",x"F7",x"BF", -- 0x4DE0
    x"FF",x"00",x"0F",x"F8",x"07",x"FF",x"DC",x"07", -- 0x4DE8
    x"FF",x"FF",x"FF",x"CF",x"FB",x"FF",x"FF",x"FF", -- 0x4DF0
    x"FF",x"FF",x"FF",x"FF",x"FC",x"00",x"00",x"00", -- 0x4DF8
    x"03",x"E0",x"0D",x"7F",x"FF",x"FF",x"F6",x"FF", -- 0x4E00
    x"FE",x"00",x"1F",x"D1",x"1F",x"FF",x"EF",x"07", -- 0x4E08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"F1",x"FF",x"FF", -- 0x4E10
    x"FF",x"FF",x"FF",x"FF",x"FE",x"00",x"00",x"00", -- 0x4E18
    x"7B",x"F0",x"0B",x"7F",x"FF",x"FF",x"F3",x"BF", -- 0x4E20
    x"FE",x"00",x"1F",x"FF",x"EF",x"FE",x"81",x"07", -- 0x4E28
    x"FF",x"FF",x"FF",x"7F",x"F8",x"40",x"FF",x"FF", -- 0x4E30
    x"FF",x"FF",x"FF",x"FF",x"FE",x"60",x"01",x"FC", -- 0x4E38
    x"1D",x"F0",x"0D",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4E40
    x"FF",x"00",x"1F",x"FF",x"01",x"FE",x"01",x"87", -- 0x4E48
    x"FE",x"EE",x"FF",x"FF",x"F0",x"00",x"1F",x"FF", -- 0x4E50
    x"FF",x"FF",x"FF",x"FF",x"FE",x"E0",x"03",x"F0", -- 0x4E58
    x"67",x"F0",x"17",x"7F",x"FF",x"FF",x"F3",x"BF", -- 0x4E60
    x"FE",x"00",x"1F",x"F8",x"01",x"FC",x"03",x"87", -- 0x4E68
    x"FF",x"FF",x"FF",x"FF",x"C0",x"00",x"0F",x"FC", -- 0x4E70
    x"3F",x"FF",x"FF",x"FF",x"FF",x"C0",x"03",x"F0", -- 0x4E78
    x"33",x"F0",x"5F",x"7F",x"FF",x"FF",x"F6",x"AF", -- 0x4E80
    x"FE",x"00",x"1F",x"FF",x"F0",x"FE",x"0F",x"87", -- 0x4E88
    x"FF",x"BF",x"FF",x"FF",x"80",x"FF",x"07",x"F8", -- 0x4E90
    x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"FA", -- 0x4E98
    x"FF",x"F1",x"BB",x"7F",x"FF",x"FF",x"F3",x"BF", -- 0x4EA0
    x"BF",x"00",x"1F",x"FF",x"FE",x"FE",x"9B",x"87", -- 0x4EA8
    x"FF",x"FF",x"FF",x"FF",x"BD",x"80",x"F3",x"F8", -- 0x4EB0
    x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"17",x"FF", -- 0x4EB8
    x"FF",x"F4",x"EE",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4EC0
    x"FF",x"00",x"1F",x"FF",x"FF",x"FF",x"03",x"87", -- 0x4EC8
    x"EF",x"EE",x"EF",x"FF",x"00",x"00",x"07",x"F8", -- 0x4ED0
    x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x4ED8
    x"FF",x"FE",x"BB",x"7F",x"FF",x"FF",x"F3",x"BF", -- 0x4EE0
    x"BF",x"00",x"0F",x"FF",x"EF",x"F8",x"83",x"87", -- 0x4EE8
    x"FF",x"FF",x"FF",x"FF",x"BE",x"BF",x"FF",x"F8", -- 0x4EF0
    x"7F",x"FF",x"FF",x"FF",x"FF",x"FD",x"B3",x"FF", -- 0x4EF8
    x"FF",x"FD",x"EE",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4F00
    x"EF",x"00",x"0F",x"FF",x"F8",x"7F",x"F7",x"8F", -- 0x4F08
    x"FF",x"FB",x"BF",x"FF",x"FF",x"FF",x"F7",x"FC", -- 0x4F10
    x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"07",x"FF", -- 0x4F18
    x"FF",x"FF",x"BB",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x4F20
    x"BB",x"00",x"0F",x"FF",x"F3",x"7F",x"0F",x"8F", -- 0x4F28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"E3",x"FC", -- 0x4F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"FF", -- 0x4F38
    x"FF",x"FF",x"EE",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4F40
    x"EF",x"00",x"0F",x"FE",x"F7",x"FF",x"CF",x"8E", -- 0x4F48
    x"FF",x"FF",x"EF",x"FF",x"FF",x"17",x"F7",x"FD", -- 0x4F50
    x"EF",x"EF",x"FE",x"FF",x"FF",x"FF",x"9F",x"FF", -- 0x4F58
    x"FF",x"FF",x"BB",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x4F60
    x"BB",x"00",x"07",x"FF",x"FE",x"FF",x"C1",x"9F", -- 0x4F68
    x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF", -- 0x4F70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"F7", -- 0x4F78
    x"FF",x"FE",x"EE",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4F80
    x"EE",x"00",x"03",x"FF",x"C4",x"1C",x"03",x"9B", -- 0x4F88
    x"FB",x"AF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x4F90
    x"FB",x"FB",x"BB",x"FF",x"BF",x"FE",x"02",x"AB", -- 0x4F98
    x"FF",x"F8",x"FB",x"7F",x"FF",x"FF",x"F3",x"BF", -- 0x4FA0
    x"BA",x"04",x"03",x"FA",x"00",x"00",x"01",x"9F", -- 0x4FA8
    x"FF",x"BB",x"FF",x"FB",x"FF",x"FF",x"FF",x"FB", -- 0x4FB0
    x"BF",x"FF",x"FB",x"FE",x"EF",x"FC",x"00",x"05", -- 0x4FB8
    x"FF",x"F9",x"EE",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x4FC0
    x"EC",x"06",x"01",x"FC",x"A2",x"00",x"03",x"9F", -- 0x4FC8
    x"EE",x"EE",x"EF",x"FE",x"FF",x"FF",x"FF",x"FE", -- 0x4FD0
    x"FF",x"FE",x"EE",x"EF",x"BF",x"FE",x"00",x"00", -- 0x4FD8
    x"3F",x"FB",x"BB",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x4FE0
    x"B0",x"00",x"01",x"FA",x"10",x"00",x"03",x"9F", -- 0x4FE8
    x"FB",x"BB",x"FF",x"FB",x"FF",x"FF",x"FF",x"FB", -- 0x4FF0
    x"BF",x"FF",x"FB",x"BE",x"EF",x"FC",x"0F",x"80", -- 0x4FF8
    x"1F",x"F6",x"EE",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x5000
    x"EE",x"00",x"00",x"68",x"5F",x"FE",x"03",x"1B", -- 0x5008
    x"AE",x"AE",x"FB",x"EE",x"FD",x"FF",x"FF",x"FE", -- 0x5010
    x"AB",x"BB",x"EA",x"FF",x"BF",x"F8",x"0B",x"FC", -- 0x5018
    x"1F",x"FF",x"BB",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x5020
    x"BA",x"00",x"00",x"7B",x"0F",x"FE",x"00",x"1F", -- 0x5028
    x"BB",x"BB",x"FF",x"FB",x"FF",x"FF",x"FF",x"FB", -- 0x5030
    x"BB",x"FF",x"BB",x"BE",x"EF",x"FC",x"07",x"FC", -- 0x5038
    x"5F",x"F6",x"EE",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x5040
    x"EE",x"00",x"00",x"14",x"40",x"3C",x"00",x"0E", -- 0x5048
    x"EE",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x5050
    x"EE",x"EE",x"EE",x"EF",x"BF",x"FE",x"00",x"61", -- 0x5058
    x"FF",x"FF",x"BB",x"7F",x"FF",x"FF",x"F3",x"BB", -- 0x5060
    x"80",x"00",x"00",x"00",x"7E",x"00",x"00",x"3F", -- 0x5068
    x"BB",x"FF",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF", -- 0x5070
    x"BB",x"FF",x"BB",x"BE",x"EF",x"FF",x"E0",x"07", -- 0x5078
    x"FF",x"FF",x"EE",x"7F",x"FF",x"FF",x"F6",x"EE", -- 0x5080
    x"00",x"00",x"00",x"00",x"3F",x"EE",x"80",x"2E", -- 0x5088
    x"AB",x"BF",x"BE",x"FC",x"FF",x"FF",x"FF",x"FE", -- 0x5090
    x"EB",x"BB",x"AA",x"BB",x"BF",x"EF",x"FA",x"FF", -- 0x5098
    x"FF",x"F8",x"0B",x"7F",x"FF",x"FF",x"F3",x"BA", -- 0x50A0
    x"00",x"00",x"C0",x"00",x"0F",x"FE",x"00",x"3B", -- 0x50A8
    x"BF",x"FF",x"FB",x"B1",x"FF",x"FF",x"FF",x"F3", -- 0x50B0
    x"BB",x"FF",x"BB",x"AE",x"EF",x"BF",x"D9",x"7F", -- 0x50B8
    x"FF",x"F8",x"02",x"7F",x"FF",x"FF",x"F6",x"EC", -- 0x50C0
    x"00",x"00",x"E0",x"00",x"00",x"00",x"00",x"EE", -- 0x50C8
    x"EE",x"EF",x"EE",x"E1",x"FF",x"FF",x"FF",x"F0", -- 0x50D0
    x"EE",x"EE",x"EE",x"EB",x"BF",x"EF",x"8E",x"3F", -- 0x50D8
    x"FF",x"F8",x"00",x"7F",x"FF",x"FF",x"F3",x"BA", -- 0x50E0
    x"00",x"00",x"F0",x"00",x"00",x"00",x"00",x"BB", -- 0x50E8
    x"BB",x"BF",x"BB",x"B1",x"FF",x"FF",x"FF",x"E0", -- 0x50F0
    x"3B",x"FF",x"BB",x"EE",x"FF",x"BB",x"00",x"5F", -- 0x50F8
    x"FF",x"F8",x"00",x"7F",x"FF",x"FF",x"F6",x"E0", -- 0x5100
    x"04",x"00",x"78",x"00",x"00",x"00",x"01",x"EE", -- 0x5108
    x"AA",x"AE",x"EA",x"C0",x"7F",x"FF",x"FF",x"80", -- 0x5110
    x"0B",x"FF",x"EF",x"AB",x"FF",x"EF",x"C2",x"3F", -- 0x5118
    x"FF",x"FF",x"E0",x"7F",x"FF",x"FF",x"F3",x"80", -- 0x5120
    x"00",x"00",x"7C",x"00",x"00",x"00",x"00",x"3B", -- 0x5128
    x"BB",x"BB",x"BB",x"00",x"3F",x"FF",x"FF",x"00", -- 0x5130
    x"03",x"FF",x"FE",x"EE",x"EF",x"BB",x"C0",x"7F", -- 0x5138
    x"FF",x"FE",x"F8",x"7F",x"FF",x"FF",x"F6",x"60", -- 0x5140
    x"C0",x"00",x"7F",x"00",x"00",x"00",x"00",x"2E", -- 0x5148
    x"EE",x"EE",x"EC",x"00",x"01",x"3F",x"FC",x"00", -- 0x5150
    x"00",x"6E",x"EF",x"FF",x"FB",x"EE",x"E2",x"3F", -- 0x5158
    x"FF",x"FE",x"78",x"7F",x"FF",x"FF",x"F0",x"98", -- 0x5160
    x"60",x"00",x"3F",x"80",x"00",x"00",x"00",x"03", -- 0x5168
    x"BB",x"BB",x"B8",x"00",x"00",x"00",x"00",x"00", -- 0x5170
    x"00",x"01",x"BB",x"BB",x"BA",x"BB",x"5F",x"9F", -- 0x5178
    x"FF",x"FC",x"F8",x"7F",x"FF",x"FF",x"F6",x"00", -- 0x5180
    x"30",x"00",x"0F",x"C0",x"00",x"00",x"00",x"00", -- 0x5188
    x"6A",x"EE",x"A0",x"00",x"00",x"00",x"00",x"00", -- 0x5190
    x"00",x"00",x"FF",x"FF",x"FA",x"EE",x"83",x"FF", -- 0x5198
    x"FF",x"FC",x"F8",x"7F",x"FF",x"FF",x"F4",x"00", -- 0x51A0
    x"00",x"00",x"07",x"E0",x"00",x"00",x"00",x"05", -- 0x51A8
    x"13",x"BB",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x51B0
    x"00",x"00",x"2E",x"EE",x"EA",x"9B",x"A3",x"FF", -- 0x51B8
    x"FF",x"FD",x"F0",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x51C0
    x"00",x"00",x"01",x"F0",x"00",x"00",x"00",x"00", -- 0x51C8
    x"0E",x"EE",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x51D0
    x"00",x"00",x"2F",x"FE",x"AA",x"0E",x"ED",x"FF", -- 0x51D8
    x"FF",x"F9",x"F0",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x51E0
    x"00",x"00",x"00",x"78",x"00",x"00",x"00",x"00", -- 0x51E8
    x"03",x"BB",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x51F0
    x"00",x"00",x"0A",x"BA",x"A8",x"0B",x"FB",x"7F", -- 0x51F8
    x"FF",x"F3",x"F0",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5200
    x"00",x"00",x"00",x"3C",x"00",x"00",x"00",x"00", -- 0x5208
    x"02",x"8A",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x5210
    x"00",x"00",x"02",x"FE",x"A0",x"06",x"FE",x"FF", -- 0x5218
    x"FF",x"07",x"F0",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5220
    x"00",x"00",x"00",x"1E",x"00",x"00",x"00",x"00", -- 0x5228
    x"07",x"03",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x5230
    x"00",x"00",x"02",x"AA",x"80",x"07",x"F9",x"FF", -- 0x5238
    x"FC",x"07",x"F4",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5240
    x"00",x"00",x"00",x"0F",x"14",x"0E",x"00",x"00", -- 0x5248
    x"02",x"80",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x5250
    x"00",x"00",x"00",x"AA",x"80",x"BF",x"FF",x"BF", -- 0x5258
    x"F0",x"0F",x"F6",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5260
    x"00",x"00",x"00",x"03",x"FF",x"FC",x"00",x"00", -- 0x5268
    x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5270
    x"00",x"00",x"00",x"EA",x"0F",x"FE",x"7C",x"77", -- 0x5278
    x"80",x"1F",x"F6",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5280
    x"00",x"00",x"00",x"01",x"FF",x"F8",x"00",x"00", -- 0x5288
    x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5290
    x"00",x"00",x"00",x"28",x"7F",x"FC",x"FE",x"80", -- 0x5298
    x"00",x"1F",x"F7",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x52A0
    x"00",x"00",x"00",x"00",x"FF",x"F0",x"00",x"00", -- 0x52A8
    x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x52B0
    x"00",x"00",x"00",x"20",x"37",x"3C",x"FE",x"C0", -- 0x52B8
    x"00",x"BF",x"F7",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x52C0
    x"00",x"00",x"00",x"07",x"7F",x"E0",x"00",x"00", -- 0x52C8
    x"F3",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x52D0
    x"00",x"00",x"00",x"00",x"3F",x"3E",x"FF",x"80", -- 0x52D8
    x"01",x"FF",x"F7",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x52E0
    x"00",x"00",x"00",x"A3",x"FF",x"C0",x"00",x"00", -- 0x52E8
    x"63",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x52F0
    x"00",x"00",x"00",x"00",x"3F",x"FD",x"EE",x"80", -- 0x52F8
    x"07",x"FF",x"F7",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5300
    x"00",x"00",x"00",x"63",x"FF",x"C0",x"00",x"00", -- 0x5308
    x"73",x"00",x"00",x"00",x"00",x"FF",x"00",x"00", -- 0x5310
    x"00",x"00",x"00",x"08",x"1F",x"78",x"F7",x"E8", -- 0x5318
    x"9F",x"FF",x"FC",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5320
    x"00",x"00",x"00",x"77",x"BF",x"80",x"00",x"00", -- 0x5328
    x"33",x"00",x"00",x"00",x"3F",x"BB",x"E0",x"00", -- 0x5330
    x"00",x"00",x"00",x"00",x"1F",x"F8",x"3B",x"55", -- 0x5338
    x"7F",x"80",x"70",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5340
    x"00",x"00",x"00",x"01",x"FF",x"00",x"00",x"00", -- 0x5348
    x"3B",x"00",x"00",x"00",x"FF",x"3B",x"FC",x"00", -- 0x5350
    x"00",x"00",x"00",x"00",x"1F",x"FF",x"1D",x"8E", -- 0x5358
    x"E7",x"82",x"F8",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5360
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00", -- 0x5368
    x"30",x"00",x"00",x"01",x"FE",x"F9",x"9F",x"00", -- 0x5370
    x"00",x"00",x"00",x"00",x"0F",x"FF",x"C1",x"17", -- 0x5378
    x"FF",x"FF",x"C0",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5380
    x"00",x"00",x"00",x"00",x"0E",x"00",x"00",x"00", -- 0x5388
    x"18",x"00",x"00",x"00",x"F8",x"FF",x"3F",x"E0", -- 0x5390
    x"00",x"04",x"00",x"00",x"0F",x"BF",x"C2",x"EF", -- 0x5398
    x"FF",x"FF",x"80",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x53A0
    x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00", -- 0x53A8
    x"1C",x"00",x"00",x"08",x"FB",x"FF",x"37",x"E0", -- 0x53B0
    x"00",x"00",x"00",x"00",x"0F",x"BF",x"C1",x"1F", -- 0x53B8
    x"FF",x"FF",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x53C0
    x"00",x"0E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x53C8
    x"0E",x"00",x"00",x"1D",x"07",x"FF",x"E3",x"68", -- 0x53D0
    x"00",x"00",x"00",x"00",x"07",x"7F",x"C7",x"3F", -- 0x53D8
    x"FF",x"FE",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x53E0
    x"00",x"00",x"00",x"00",x"1C",x"00",x"00",x"00", -- 0x53E8
    x"00",x"00",x"00",x"00",x"3F",x"FF",x"FB",x"F6", -- 0x53F0
    x"00",x"00",x"00",x"00",x"07",x"7F",x"E1",x"7F", -- 0x53F8
    x"FF",x"FC",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5400
    x"00",x"00",x"00",x"00",x"0E",x"00",x"00",x"00", -- 0x5408
    x"00",x"00",x"01",x"C6",x"7F",x"FF",x"FF",x"E8", -- 0x5410
    x"00",x"00",x"00",x"00",x"07",x"0F",x"F3",x"8F", -- 0x5418
    x"97",x"FC",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5420
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5428
    x"00",x"00",x"01",x"B1",x"EF",x"FF",x"EF",x"B7", -- 0x5430
    x"00",x"00",x"00",x"00",x"07",x"83",x"E1",x"C6", -- 0x5438
    x"00",x"78",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5440
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5448
    x"00",x"00",x"00",x"21",x"DF",x"FF",x"D1",x"A2", -- 0x5450
    x"00",x"00",x"40",x"00",x"03",x"00",x"F1",x"FF", -- 0x5458
    x"14",x"20",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5460
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5468
    x"00",x"00",x"00",x"3E",x"FF",x"FF",x"FF",x"DF", -- 0x5470
    x"00",x"00",x"00",x"00",x"03",x"06",x"70",x"7C", -- 0x5478
    x"00",x"C0",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5480
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5488
    x"00",x"00",x"00",x"0F",x"FF",x"FF",x"FF",x"E7", -- 0x5490
    x"E0",x"00",x"00",x"00",x"03",x"87",x"F1",x"F8", -- 0x5498
    x"03",x"80",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x54A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x54A8
    x"00",x"00",x"00",x"1E",x"AF",x"FF",x"FF",x"F7", -- 0x54B0
    x"00",x"00",x"00",x"00",x"03",x"8F",x"FB",x"F8", -- 0x54B8
    x"20",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x54C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x54C8
    x"00",x"00",x"00",x"1F",x"BF",x"FF",x"FF",x"BF", -- 0x54D0
    x"E0",x"00",x"00",x"00",x"F3",x"8D",x"FF",x"F8", -- 0x54D8
    x"5F",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x54E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x54E8
    x"00",x"00",x"00",x"1E",x"FF",x"FF",x"FF",x"4F", -- 0x54F0
    x"F0",x"00",x"00",x"01",x"E3",x"87",x"FF",x"FC", -- 0x54F8
    x"6E",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5500
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5508
    x"00",x"00",x"00",x"0D",x"F7",x"BF",x"FF",x"EF", -- 0x5510
    x"E8",x"00",x"00",x"00",x"01",x"1F",x"FF",x"FF", -- 0x5518
    x"FE",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5520
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5528
    x"00",x"00",x"00",x"0B",x"FF",x"9F",x"FF",x"FD", -- 0x5530
    x"F8",x"00",x"00",x"00",x"01",x"BF",x"FF",x"FF", -- 0x5538
    x"FF",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5540
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5548
    x"00",x"00",x"00",x"07",x"FF",x"FF",x"FF",x"8F", -- 0x5550
    x"E8",x"00",x"00",x"00",x"01",x"BF",x"FF",x"FF", -- 0x5558
    x"FC",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5560
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5568
    x"00",x"00",x"00",x"07",x"FF",x"FF",x"FF",x"FF", -- 0x5570
    x"F8",x"00",x"00",x"00",x"01",x"BF",x"FF",x"FF", -- 0x5578
    x"F8",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5580
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5588
    x"00",x"00",x"00",x"07",x"FF",x"FF",x"9F",x"FF", -- 0x5590
    x"F8",x"00",x"00",x"00",x"01",x"3F",x"FF",x"FF", -- 0x5598
    x"F0",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x55A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x55A8
    x"FE",x"00",x"00",x"07",x"FF",x"1F",x"FF",x"F5", -- 0x55B0
    x"FC",x"00",x"00",x"00",x"01",x"3F",x"FF",x"FF", -- 0x55B8
    x"E0",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x55C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x55C8
    x"00",x"00",x"00",x"03",x"FC",x"3F",x"FF",x"BF", -- 0x55D0
    x"F8",x"00",x"00",x"00",x"01",x"3F",x"85",x"FF", -- 0x55D8
    x"C0",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x55E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x55E8
    x"00",x"00",x"00",x"03",x"FF",x"F7",x"FF",x"DF", -- 0x55F0
    x"F8",x"00",x"00",x"00",x"00",x"1D",x"2A",x"07", -- 0x55F8
    x"80",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5600
    x"00",x"0E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5608
    x"00",x"00",x"00",x"07",x"FF",x"FF",x"FF",x"FF", -- 0x5610
    x"F8",x"00",x"00",x"00",x"01",x"06",x"FF",x"00", -- 0x5618
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5620
    x"00",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5628
    x"10",x"00",x"00",x"1F",x"FF",x"FF",x"FF",x"DF", -- 0x5630
    x"F8",x"00",x"00",x"00",x"01",x"17",x"3D",x"95", -- 0x5638
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5640
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01", -- 0x5648
    x"FF",x"80",x"00",x"07",x"FF",x"FF",x"FF",x"EF", -- 0x5650
    x"F8",x"00",x"00",x"00",x"00",x"0E",x"EF",x"DA", -- 0x5658
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5660
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5668
    x"00",x"00",x"00",x"03",x"FF",x"FF",x"FF",x"F7", -- 0x5670
    x"F0",x"00",x"00",x"00",x"00",x"15",x"F7",x"80", -- 0x5678
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5680
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5688
    x"00",x"00",x"00",x"03",x"FF",x"FF",x"FF",x"ED", -- 0x5690
    x"E0",x"00",x"00",x"00",x"00",x"0F",x"BF",x"EC", -- 0x5698
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x56A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x56A8
    x"00",x"00",x"00",x"07",x"FF",x"FF",x"FF",x"DC", -- 0x56B0
    x"E0",x"00",x"00",x"00",x"00",x"17",x"7F",x"D8", -- 0x56B8
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x56C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x56C8
    x"00",x"00",x"00",x"07",x"FF",x"FF",x"FF",x"BC", -- 0x56D0
    x"C0",x"00",x"00",x"00",x"00",x"3F",x"FF",x"F8", -- 0x56D8
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x56E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x56E8
    x"00",x"00",x"00",x"03",x"FF",x"FF",x"FF",x"DE", -- 0x56F0
    x"00",x"00",x"00",x"00",x"00",x"7F",x"FF",x"F8", -- 0x56F8
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5700
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5708
    x"00",x"00",x"00",x"01",x"FF",x"FF",x"FF",x"FF", -- 0x5710
    x"80",x"00",x"00",x"00",x"00",x"7F",x"FF",x"F8", -- 0x5718
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5720
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5728
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"FF", -- 0x5730
    x"80",x"00",x"00",x"00",x"00",x"7F",x"FF",x"F0", -- 0x5738
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5740
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5748
    x"00",x"00",x"00",x"03",x"DF",x"FE",x"C1",x"F2", -- 0x5750
    x"00",x"00",x"00",x"00",x"18",x"7F",x"FF",x"F0", -- 0x5758
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5760
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5768
    x"00",x"00",x"00",x"00",x"83",x"00",x"1F",x"CC", -- 0x5770
    x"00",x"00",x"00",x"00",x"00",x"7F",x"FF",x"F0", -- 0x5778
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5780
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5788
    x"00",x"00",x"00",x"03",x"00",x"80",x"3F",x"98", -- 0x5790
    x"00",x"00",x"00",x"00",x"00",x"7F",x"FF",x"F0", -- 0x5798
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x57A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x57A8
    x"00",x"00",x"00",x"00",x"E2",x"46",x"3E",x"60", -- 0x57B0
    x"00",x"00",x"00",x"00",x"00",x"7F",x"FF",x"E0", -- 0x57B8
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x57C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x57C8
    x"00",x"00",x"00",x"01",x"80",x"33",x"3C",x"00", -- 0x57D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"60", -- 0x57D8
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x57E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x57E8
    x"00",x"00",x"00",x"00",x"A0",x"73",x"10",x"00", -- 0x57F0
    x"00",x"00",x"00",x"00",x"00",x"15",x"3A",x"80", -- 0x57F8
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5800
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5808
    x"00",x"00",x"00",x"00",x"E0",x"08",x"18",x"00", -- 0x5810
    x"00",x"00",x"00",x"00",x"00",x"02",x"F6",x"00", -- 0x5818
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5820
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5828
    x"00",x"00",x"00",x"00",x"E0",x"00",x"00",x"00", -- 0x5830
    x"00",x"00",x"00",x"00",x"00",x"17",x"B6",x"00", -- 0x5838
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5840
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5848
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5850
    x"00",x"00",x"00",x"00",x"00",x"02",x"ED",x"80", -- 0x5858
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5860
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5868
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5870
    x"00",x"00",x"00",x"00",x"00",x"05",x"2C",x"00", -- 0x5878
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5880
    x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5888
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5890
    x"00",x"00",x"00",x"00",x"00",x"02",x"B0",x"80", -- 0x5898
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x58A0
    x"00",x"70",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x58A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x58B0
    x"00",x"00",x"00",x"00",x"00",x"7F",x"FF",x"00", -- 0x58B8
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x58C0
    x"00",x"78",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x58C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x58D0
    x"00",x"40",x"00",x"00",x"00",x"7F",x"FF",x"80", -- 0x58D8
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x58E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x58E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x58F0
    x"00",x"40",x"00",x"00",x"00",x"7F",x"FF",x"C0", -- 0x58F8
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5900
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5908
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5910
    x"00",x"00",x"00",x"00",x"00",x"7F",x"FF",x"80", -- 0x5918
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5920
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5928
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5930
    x"00",x"00",x"00",x"00",x"00",x"7F",x"FF",x"80", -- 0x5938
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5940
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5948
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5950
    x"00",x"00",x"00",x"00",x"00",x"7F",x"FF",x"80", -- 0x5958
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5960
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5968
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5970
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5978
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5980
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5988
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5990
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5998
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x59A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x59A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x59B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x59B8
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x59C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x59C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x59D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x59D8
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x59E0
    x"FF",x"3C",x"FF",x"F3",x"3F",x"FF",x"CF",x"9F", -- 0x59E8
    x"FF",x"FF",x"FF",x"03",x"FF",x"CC",x"FF",x"FF", -- 0x59F0
    x"F3",x"FF",x"FF",x"F8",x"1F",x"FE",x"0F",x"FF", -- 0x59F8
    x"8F",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5A00
    x"FF",x"18",x"FF",x"F3",x"3F",x"FF",x"CF",x"FF", -- 0x5A08
    x"FF",x"FF",x"FF",x"CF",x"FF",x"CC",x"FF",x"FF", -- 0x5A10
    x"FF",x"FF",x"FF",x"FE",x"7F",x"FE",x"7F",x"FF", -- 0x5A18
    x"CF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5A20
    x"FF",x"00",x"FF",x"F3",x"31",x"9E",x"49",x"10", -- 0x5A28
    x"E1",x"FF",x"FF",x"CF",x"FF",x"CC",x"C6",x"08", -- 0x5A30
    x"23",x"0F",x"FF",x"FE",x"7F",x"FE",x"7C",x"60", -- 0x5A38
    x"CC",x"70",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5A40
    x"FF",x"24",x"FF",x"F0",x"3C",x"C0",x"C3",x"92", -- 0x5A48
    x"4F",x"FF",x"FF",x"CF",x"FF",x"C0",x"F2",x"38", -- 0x5A50
    x"F2",x"7F",x"FF",x"FE",x"7F",x"FE",x"1F",x"23", -- 0x5A58
    x"C9",x"27",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5A60
    x"FF",x"3C",x"FF",x"F3",x"30",x"C0",x"C7",x"92", -- 0x5A68
    x"63",x"FF",x"FF",x"CF",x"FF",x"CC",x"C2",x"79", -- 0x5A70
    x"F3",x"1F",x"FF",x"FE",x"7F",x"FE",x"7C",x"27", -- 0x5A78
    x"C8",x"31",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5A80
    x"FF",x"3C",x"FF",x"F3",x"24",x"E1",x"C3",x"92", -- 0x5A88
    x"79",x"FF",x"FF",x"CF",x"FF",x"CC",x"92",x"79", -- 0x5A90
    x"F3",x"CF",x"FF",x"FE",x"7F",x"FE",x"79",x"27", -- 0x5A98
    x"C9",x"FC",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5AA0
    x"FF",x"3C",x"9F",x"F3",x"30",x"E1",x"C9",x"92", -- 0x5AA8
    x"43",x"FF",x"FF",x"CE",x"7F",x"CC",x"C2",x"79", -- 0x5AB0
    x"F2",x"1F",x"FF",x"FE",x"73",x"FE",x"0C",x"27", -- 0x5AB8
    x"CC",x"61",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5AC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5AC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5AD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5AD8
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5AE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5AE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5AF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5AF8
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5B00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B18
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5B20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B38
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F7",x"FF", -- 0x5B40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B58
    x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"F0",x"00", -- 0x5B60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5B70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5B78
    x"00",x"00",x"00",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x5B80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5B98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5BF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00", -- 0x5C00
    x"A0",x"27",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5C08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5C10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5C18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5C20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5C28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5C30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5C38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5C40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5C48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5C50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5C58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5C68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5C78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5C88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5C98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5CA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5CB8
    x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5CC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5CD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5CE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5CF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5D00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5D08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5D10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5D20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5D28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5D30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5D38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5D40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5D48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5D50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5D60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5D68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5D70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5D80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5D88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5D90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5DA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5DA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5DB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5DB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5DC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5DC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5DD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5DD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5DE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5DF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5DF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5E08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5E18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5E28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5E38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5E48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5E58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5E68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5E78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5E88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5E98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5EA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5EB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5EC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5ED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5EE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5F00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5F10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5F20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5F40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5F50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5F60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5F70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5F80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5F90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5FA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5FB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5FC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5FC8
    x"00",x"00",x"00",x"40",x"00",x"00",x"00",x"00", -- 0x5FD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5FE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x5FF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x5FF8
    x"00",x"E6",x"E0",x"19",x"E0",x"4D",x"E0",x"97", -- 0x6000
    x"E0",x"B5",x"E0",x"A1",x"E0",x"FF",x"E1",x"19", -- 0x6008
    x"7E",x"A0",x"5E",x"00",x"00",x"00",x"00",x"00", -- 0x6010
    x"00",x"34",x"32",x"10",x"21",x"1F",x"E1",x"8E", -- 0x6018
    x"E0",x"32",x"96",x"E7",x"27",x"5C",x"8E",x"E0", -- 0x6020
    x"3B",x"81",x"01",x"27",x"55",x"8E",x"E0",x"44", -- 0x6028
    x"20",x"50",x"CC",x"00",x"00",x"00",x"00",x"0F", -- 0x6030
    x"E0",x"00",x"00",x"4C",x"03",x"05",x"12",x"00", -- 0x6038
    x"00",x"D8",x"00",x"00",x"4C",x"03",x"15",x"12", -- 0x6040
    x"00",x"00",x"D8",x"00",x"00",x"34",x"32",x"10", -- 0x6048
    x"21",x"1F",x"AD",x"8E",x"E0",x"70",x"10",x"8E", -- 0x6050
    x"E0",x"6C",x"96",x"E6",x"81",x"02",x"23",x"03", -- 0x6058
    x"8E",x"E0",x"79",x"80",x"01",x"A6",x"A6",x"A7", -- 0x6060
    x"02",x"7E",x"E0",x"82",x"15",x"1E",x"14",x"1D", -- 0x6068
    x"4C",x"80",x"00",x"00",x"00",x"00",x"C0",x"00", -- 0x6070
    x"00",x"4C",x"80",x"00",x"00",x"00",x"00",x"C0", -- 0x6078
    x"00",x"00",x"A6",x"80",x"B7",x"FF",x"90",x"10", -- 0x6080
    x"8E",x"FF",x"98",x"A6",x"80",x"A7",x"A0",x"10", -- 0x6088
    x"8C",x"FF",x"A0",x"25",x"F6",x"35",x"B2",x"34", -- 0x6090
    x"36",x"30",x"8D",x"00",x"44",x"8D",x"52",x"35", -- 0x6098
    x"B6",x"34",x"36",x"30",x"8D",x"00",x"3A",x"34", -- 0x60A0
    x"10",x"E7",x"84",x"8D",x"44",x"C6",x"38",x"35", -- 0x60A8
    x"10",x"E7",x"84",x"35",x"B6",x"34",x"36",x"30", -- 0x60B0
    x"8D",x"00",x"26",x"34",x"10",x"C6",x"36",x"E7", -- 0x60B8
    x"01",x"8D",x"2E",x"35",x"10",x"C6",x"39",x"E7", -- 0x60C0
    x"01",x"35",x"B6",x"34",x"36",x"30",x"8D",x"00", -- 0x60C8
    x"10",x"34",x"10",x"C6",x"34",x"E7",x"0E",x"8D", -- 0x60D0
    x"18",x"35",x"10",x"C6",x"35",x"E7",x"0E",x"35", -- 0x60D8
    x"B6",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E", -- 0x60E0
    x"3F",x"38",x"30",x"31",x"32",x"33",x"3D",x"35", -- 0x60E8
    x"3F",x"10",x"8E",x"FF",x"A0",x"C6",x"10",x"A6", -- 0x60F0
    x"80",x"A7",x"A0",x"5A",x"26",x"F9",x"39",x"DD", -- 0x60F8
    x"40",x"EC",x"E4",x"DD",x"42",x"EC",x"62",x"DD", -- 0x6100
    x"44",x"5F",x"F7",x"FF",x"91",x"10",x"DE",x"44", -- 0x6108
    x"DC",x"42",x"34",x"06",x"DC",x"40",x"1C",x"AF", -- 0x6110
    x"39",x"1A",x"50",x"DD",x"40",x"35",x"06",x"DD", -- 0x6118
    x"42",x"10",x"DF",x"44",x"C6",x"01",x"F7",x"FF", -- 0x6120
    x"91",x"10",x"CE",x"DF",x"FF",x"DC",x"44",x"34", -- 0x6128
    x"06",x"DC",x"42",x"34",x"06",x"DC",x"40",x"39", -- 0x6130
    x"0D",x"41",x"26",x"16",x"96",x"42",x"81",x"62", -- 0x6138
    x"23",x"06",x"CE",x"01",x"1B",x"7E",x"B8",x"D7", -- 0x6140
    x"86",x"62",x"CE",x"E1",x"58",x"97",x"42",x"7E", -- 0x6148
    x"B8",x"9D",x"96",x"42",x"81",x"29",x"23",x"03", -- 0x6150
    x"7E",x"B8",x"D7",x"86",x"29",x"CE",x"E1",x"5D", -- 0x6158
    x"20",x"EB",x"17",x"E1",x"C5",x"E1",x"92",x"05", -- 0x6160
    x"E2",x"64",x"E1",x"A6",x"00",x"00",x"00",x"00", -- 0x6168
    x"00",x"00",x"33",x"4A",x"6D",x"C4",x"10",x"26", -- 0x6170
    x"D6",x"7F",x"30",x"1F",x"A6",x"80",x"84",x"7F", -- 0x6178
    x"81",x"62",x"25",x"07",x"80",x"62",x"CE",x"E1", -- 0x6180
    x"58",x"20",x"E7",x"80",x"29",x"CE",x"E1",x"5D", -- 0x6188
    x"20",x"E0",x"81",x"E2",x"25",x"04",x"81",x"F8", -- 0x6190
    x"23",x"04",x"6E",x"9F",x"01",x"37",x"80",x"E2", -- 0x6198
    x"8E",x"E2",x"36",x"7E",x"AD",x"D4",x"C1",x"52", -- 0x61A0
    x"25",x"04",x"C1",x"5A",x"23",x"04",x"6E",x"9F", -- 0x61A8
    x"01",x"3C",x"C0",x"52",x"C1",x"04",x"24",x"07", -- 0x61B0
    x"34",x"04",x"BD",x"B2",x"62",x"35",x"04",x"8E", -- 0x61B8
    x"E2",x"7E",x"7E",x"B2",x"CE",x"57",x"49",x"44", -- 0x61C0
    x"54",x"C8",x"50",x"41",x"4C",x"45",x"54",x"54", -- 0x61C8
    x"C5",x"48",x"53",x"43",x"52",x"45",x"45",x"CE", -- 0x61D0
    x"4C",x"50",x"4F",x"4B",x"C5",x"48",x"43",x"4C", -- 0x61D8
    x"D3",x"48",x"43",x"4F",x"4C",x"4F",x"D2",x"48", -- 0x61E0
    x"50",x"41",x"49",x"4E",x"D4",x"48",x"43",x"49", -- 0x61E8
    x"52",x"43",x"4C",x"C5",x"48",x"4C",x"49",x"4E", -- 0x61F0
    x"C5",x"48",x"47",x"45",x"D4",x"48",x"50",x"55", -- 0x61F8
    x"D4",x"48",x"42",x"55",x"46",x"C6",x"48",x"50", -- 0x6200
    x"52",x"49",x"4E",x"D4",x"45",x"52",x"D2",x"42", -- 0x6208
    x"52",x"CB",x"4C",x"4F",x"43",x"41",x"54",x"C5", -- 0x6210
    x"48",x"53",x"54",x"41",x"D4",x"48",x"53",x"45", -- 0x6218
    x"D4",x"48",x"52",x"45",x"53",x"45",x"D4",x"48", -- 0x6220
    x"44",x"52",x"41",x"D7",x"43",x"4D",x"D0",x"52", -- 0x6228
    x"47",x"C2",x"41",x"54",x"54",x"D2",x"F6",x"36", -- 0x6230
    x"E5",x"F0",x"E6",x"88",x"E5",x"45",x"E6",x"CF", -- 0x6238
    x"E6",x"F4",x"EB",x"F5",x"EA",x"49",x"E8",x"82", -- 0x6240
    x"ED",x"E5",x"ED",x"ED",x"ED",x"58",x"EF",x"3F", -- 0x6248
    x"E3",x"D4",x"E3",x"E6",x"F8",x"D2",x"F9",x"25", -- 0x6250
    x"E7",x"61",x"E7",x"65",x"F3",x"9D",x"E6",x"76", -- 0x6258
    x"E6",x"74",x"F9",x"B9",x"4C",x"50",x"45",x"45", -- 0x6260
    x"CB",x"42",x"55",x"54",x"54",x"4F",x"CE",x"48", -- 0x6268
    x"50",x"4F",x"49",x"4E",x"D4",x"45",x"52",x"4E", -- 0x6270
    x"CF",x"45",x"52",x"4C",x"49",x"CE",x"E5",x"73", -- 0x6278
    x"E5",x"B1",x"E8",x"5C",x"E4",x"E9",x"E4",x"FD", -- 0x6280
    x"8E",x"80",x"E7",x"BD",x"B9",x"9C",x"8E",x"E2", -- 0x6288
    x"F7",x"BD",x"B9",x"9C",x"7E",x"80",x"B8",x"8E", -- 0x6290
    x"E2",x"A2",x"7E",x"C0",x"C9",x"8E",x"E3",x"15", -- 0x6298
    x"7E",x"C0",x"DC",x"44",x"49",x"53",x"4B",x"20", -- 0x62A0
    x"45",x"58",x"54",x"45",x"4E",x"44",x"45",x"44", -- 0x62A8
    x"20",x"43",x"4F",x"4C",x"4F",x"52",x"20",x"42", -- 0x62B0
    x"41",x"53",x"49",x"43",x"20",x"32",x"2E",x"30", -- 0x62B8
    x"0D",x"43",x"4F",x"50",x"52",x"2E",x"20",x"31", -- 0x62C0
    x"39",x"38",x"31",x"2C",x"20",x"31",x"39",x"38", -- 0x62C8
    x"36",x"20",x"42",x"59",x"20",x"54",x"41",x"4E", -- 0x62D0
    x"44",x"59",x"0D",x"55",x"4E",x"44",x"45",x"52", -- 0x62D8
    x"20",x"4C",x"49",x"43",x"45",x"4E",x"53",x"45", -- 0x62E0
    x"20",x"46",x"52",x"4F",x"4D",x"20",x"4D",x"49", -- 0x62E8
    x"43",x"52",x"4F",x"53",x"4F",x"46",x"54",x"0D", -- 0x62F0
    x"41",x"4E",x"44",x"20",x"4D",x"49",x"43",x"52", -- 0x62F8
    x"4F",x"57",x"41",x"52",x"45",x"20",x"53",x"59", -- 0x6300
    x"53",x"54",x"45",x"4D",x"53",x"20",x"43",x"4F", -- 0x6308
    x"52",x"50",x"2E",x"0D",x"0D",x"00",x"44",x"49", -- 0x6310
    x"53",x"4B",x"20",x"45",x"58",x"54",x"45",x"4E", -- 0x6318
    x"44",x"45",x"44",x"20",x"43",x"4F",x"4C",x"4F", -- 0x6320
    x"52",x"20",x"42",x"41",x"53",x"49",x"43",x"20", -- 0x6328
    x"32",x"2E",x"31",x"0D",x"43",x"4F",x"50",x"52", -- 0x6330
    x"2E",x"20",x"31",x"39",x"38",x"32",x"2C",x"20", -- 0x6338
    x"31",x"39",x"38",x"36",x"20",x"42",x"59",x"20", -- 0x6340
    x"54",x"41",x"4E",x"44",x"59",x"0D",x"55",x"4E", -- 0x6348
    x"44",x"45",x"52",x"20",x"4C",x"49",x"43",x"45", -- 0x6350
    x"4E",x"53",x"45",x"20",x"46",x"52",x"4F",x"4D", -- 0x6358
    x"20",x"4D",x"49",x"43",x"52",x"4F",x"53",x"4F", -- 0x6360
    x"46",x"54",x"0D",x"41",x"4E",x"44",x"20",x"4D", -- 0x6368
    x"49",x"43",x"52",x"4F",x"57",x"41",x"52",x"45", -- 0x6370
    x"20",x"53",x"59",x"53",x"54",x"45",x"4D",x"53", -- 0x6378
    x"20",x"43",x"4F",x"52",x"50",x"2E",x"0D",x"0D", -- 0x6380
    x"00",x"4F",x"5F",x"10",x"21",x"1C",x"71",x"F7", -- 0x6388
    x"FE",x"08",x"DD",x"E6",x"FD",x"FE",x"0C",x"FD", -- 0x6390
    x"FE",x"0E",x"B7",x"FE",x"0B",x"86",x"01",x"B7", -- 0x6398
    x"FE",x"0A",x"86",x"34",x"B7",x"FF",x"A0",x"CC", -- 0x63A0
    x"FF",x"FF",x"DD",x"00",x"86",x"38",x"B7",x"FF", -- 0x63A8
    x"A0",x"7E",x"AD",x"19",x"81",x"EF",x"27",x"1C", -- 0x63B0
    x"81",x"F0",x"27",x"2A",x"BD",x"B7",x"0B",x"7E", -- 0x63B8
    x"AF",x"45",x"9D",x"9F",x"81",x"81",x"26",x"07", -- 0x63C0
    x"9D",x"9F",x"81",x"A5",x"26",x"01",x"39",x"32", -- 0x63C8
    x"62",x"7E",x"B2",x"77",x"8D",x"EC",x"9D",x"9F", -- 0x63D0
    x"BD",x"AF",x"67",x"DC",x"2B",x"FD",x"FE",x"0E", -- 0x63D8
    x"DC",x"68",x"FD",x"FE",x"11",x"39",x"8D",x"DA", -- 0x63E0
    x"9D",x"9F",x"BD",x"AF",x"67",x"DC",x"2B",x"FD", -- 0x63E8
    x"FE",x"0C",x"DC",x"68",x"FD",x"FE",x"15",x"39", -- 0x63F0
    x"68",x"02",x"69",x"01",x"69",x"84",x"10",x"25", -- 0x63F8
    x"D6",x"90",x"5A",x"26",x"F3",x"80",x"30",x"AB", -- 0x6400
    x"02",x"A7",x"02",x"39",x"10",x"25",x"A3",x"F0", -- 0x6408
    x"7E",x"88",x"3F",x"81",x"03",x"1A",x"01",x"26", -- 0x6410
    x"0D",x"34",x"03",x"96",x"E6",x"27",x"05",x"0F", -- 0x6418
    x"E6",x"BD",x"E0",x"19",x"35",x"03",x"7E",x"A3", -- 0x6420
    x"C6",x"81",x"03",x"27",x"03",x"7E",x"AD",x"F4", -- 0x6428
    x"86",x"01",x"B7",x"FE",x"17",x"96",x"68",x"4C", -- 0x6430
    x"27",x"05",x"FC",x"FE",x"0C",x"26",x"0A",x"96", -- 0x6438
    x"E6",x"27",x"03",x"BD",x"E0",x"19",x"7E",x"AE", -- 0x6440
    x"09",x"DD",x"2B",x"7D",x"FE",x"17",x"26",x"08", -- 0x6448
    x"10",x"DE",x"21",x"CC",x"AD",x"C4",x"34",x"06", -- 0x6450
    x"BD",x"AE",x"EB",x"30",x"01",x"DC",x"2B",x"10", -- 0x6458
    x"93",x"68",x"22",x"02",x"9E",x"19",x"BD",x"AD", -- 0x6460
    x"05",x"10",x"25",x"00",x"B1",x"7E",x"AE",x"BB", -- 0x6468
    x"7F",x"FE",x"17",x"96",x"68",x"4C",x"27",x"05", -- 0x6470
    x"BE",x"FE",x"0E",x"26",x"36",x"34",x"02",x"96", -- 0x6478
    x"E6",x"35",x"02",x"27",x"03",x"BD",x"E0",x"19", -- 0x6480
    x"C1",x"4C",x"26",x"13",x"BD",x"B9",x"5C",x"BD", -- 0x6488
    x"B9",x"AF",x"30",x"8D",x"00",x"36",x"BD",x"AC", -- 0x6490
    x"A0",x"BD",x"AC",x"A0",x"7E",x"AC",x"65",x"C1", -- 0x6498
    x"4E",x"26",x"0D",x"BD",x"B9",x"5C",x"BD",x"B9", -- 0x64A0
    x"AF",x"30",x"8D",x"00",x"21",x"7E",x"E4",x"96", -- 0x64A8
    x"7E",x"AC",x"49",x"F7",x"FE",x"10",x"34",x"04", -- 0x64B0
    x"DC",x"68",x"FD",x"FE",x"13",x"35",x"04",x"C1", -- 0x64B8
    x"06",x"26",x"04",x"DC",x"2B",x"DD",x"A6",x"1F", -- 0x64C0
    x"10",x"16",x"FF",x"7D",x"48",x"52",x"48",x"50", -- 0x64C8
    x"34",x"06",x"4F",x"5F",x"DD",x"2D",x"FD",x"FE", -- 0x64D0
    x"0C",x"FD",x"FE",x"0E",x"FD",x"FE",x"13",x"86", -- 0x64D8
    x"FF",x"B7",x"FE",x"10",x"35",x"06",x"7E",x"AD", -- 0x64E0
    x"43",x"4F",x"F6",x"FE",x"10",x"C1",x"FF",x"26", -- 0x64E8
    x"03",x"1D",x"20",x"06",x"C1",x"F1",x"26",x"01", -- 0x64F0
    x"53",x"57",x"7E",x"B4",x"F4",x"FC",x"FE",x"13", -- 0x64F8
    x"20",x"F8",x"BD",x"E0",x"19",x"BD",x"B9",x"5C", -- 0x6500
    x"1A",x"50",x"86",x"34",x"B7",x"FF",x"A0",x"CC", -- 0x6508
    x"FF",x"FF",x"DD",x"00",x"86",x"38",x"B7",x"FF", -- 0x6510
    x"A0",x"1C",x"AF",x"7E",x"AC",x"76",x"7D",x"FE", -- 0x6518
    x"17",x"27",x"05",x"FC",x"FE",x"15",x"20",x"03", -- 0x6520
    x"FC",x"FE",x"11",x"DD",x"68",x"C6",x"0E",x"7E", -- 0x6528
    x"AC",x"49",x"FC",x"FE",x"0C",x"10",x"27",x"C8", -- 0x6530
    x"D8",x"34",x"06",x"86",x"01",x"B7",x"FE",x"17", -- 0x6538
    x"35",x"06",x"16",x"FF",x"04",x"BD",x"B1",x"41", -- 0x6540
    x"10",x"21",x"1A",x"B4",x"8D",x"40",x"C1",x"3F", -- 0x6548
    x"10",x"22",x"CE",x"F6",x"34",x"14",x"BD",x"B2", -- 0x6550
    x"6D",x"BD",x"B7",x"0B",x"1F",x"98",x"35",x"14", -- 0x6558
    x"C1",x"3F",x"10",x"22",x"CE",x"E4",x"1A",x"50", -- 0x6560
    x"17",x"FB",x"36",x"A7",x"84",x"17",x"FB",x"27", -- 0x6568
    x"1C",x"AF",x"39",x"8D",x"19",x"10",x"21",x"1A", -- 0x6570
    x"87",x"C1",x"3F",x"10",x"22",x"CE",x"CB",x"1A", -- 0x6578
    x"50",x"17",x"FB",x"1D",x"E6",x"84",x"17",x"FB", -- 0x6580
    x"0E",x"1C",x"AF",x"7E",x"B4",x"F3",x"34",x"02", -- 0x6588
    x"96",x"4F",x"81",x"93",x"23",x"04",x"C6",x"40", -- 0x6590
    x"20",x"15",x"BD",x"BC",x"C8",x"DC",x"52",x"84", -- 0x6598
    x"1F",x"1F",x"01",x"DC",x"51",x"47",x"56",x"47", -- 0x65A0
    x"56",x"47",x"56",x"47",x"56",x"47",x"56",x"35", -- 0x65A8
    x"82",x"BD",x"B3",x"ED",x"10",x"21",x"1A",x"48", -- 0x65B0
    x"C1",x"03",x"10",x"22",x"CE",x"8C",x"1F",x"98", -- 0x65B8
    x"5F",x"53",x"8E",x"FF",x"00",x"E7",x"02",x"E6", -- 0x65C0
    x"84",x"C1",x"0F",x"27",x"1D",x"30",x"8D",x"00", -- 0x65C8
    x"04",x"48",x"48",x"6E",x"86",x"C4",x"01",x"20", -- 0x65D0
    x"0A",x"C4",x"04",x"20",x"06",x"C4",x"02",x"20", -- 0x65D8
    x"02",x"C4",x"08",x"26",x"05",x"CC",x"00",x"01", -- 0x65E0
    x"20",x"02",x"4F",x"5F",x"BD",x"B4",x"F4",x"39", -- 0x65E8
    x"81",x"F7",x"10",x"21",x"1A",x"0A",x"26",x"08", -- 0x65F0
    x"9D",x"9F",x"30",x"8D",x"00",x"66",x"20",x"34", -- 0x65F8
    x"81",x"F6",x"26",x"08",x"9D",x"9F",x"30",x"8D", -- 0x6600
    x"00",x"4A",x"20",x"28",x"BD",x"E7",x"B2",x"8E", -- 0x6608
    x"FF",x"B0",x"10",x"8E",x"E6",x"78",x"96",x"2C", -- 0x6610
    x"81",x"10",x"10",x"24",x"CE",x"2C",x"30",x"86", -- 0x6618
    x"31",x"A6",x"D6",x"C0",x"C1",x"3F",x"23",x"02", -- 0x6620
    x"C6",x"3F",x"1A",x"50",x"13",x"E7",x"84",x"E7", -- 0x6628
    x"A4",x"1C",x"AF",x"39",x"34",x"10",x"10",x"8E", -- 0x6630
    x"E6",x"78",x"8D",x"0C",x"35",x"10",x"10",x"8E", -- 0x6638
    x"FF",x"B0",x"1A",x"50",x"13",x"8D",x"01",x"39", -- 0x6640
    x"C6",x"0F",x"A6",x"80",x"A7",x"A0",x"5A",x"26", -- 0x6648
    x"F9",x"1C",x"AF",x"39",x"12",x"24",x"0B",x"07", -- 0x6650
    x"3F",x"1F",x"09",x"26",x"00",x"12",x"00",x"3F", -- 0x6658
    x"00",x"12",x"00",x"26",x"12",x"36",x"09",x"24", -- 0x6660
    x"3F",x"1B",x"2D",x"26",x"00",x"12",x"00",x"3F", -- 0x6668
    x"00",x"12",x"00",x"26",x"20",x"84",x"20",x"8E", -- 0x6670
    x"12",x"24",x"0B",x"07",x"3F",x"1F",x"09",x"26", -- 0x6678
    x"00",x"12",x"00",x"3F",x"00",x"12",x"00",x"26", -- 0x6680
    x"81",x"00",x"10",x"21",x"19",x"72",x"26",x"03", -- 0x6688
    x"5F",x"20",x"09",x"BD",x"B7",x"0B",x"C1",x"04", -- 0x6690
    x"10",x"22",x"CD",x"AE",x"D7",x"E6",x"C1",x"00", -- 0x6698
    x"26",x"03",x"7E",x"E0",x"19",x"D7",x"E6",x"8E", -- 0x66A0
    x"E6",x"CB",x"C0",x"01",x"A6",x"85",x"97",x"B9", -- 0x66A8
    x"C1",x"01",x"2E",x"05",x"CC",x"00",x"A0",x"20", -- 0x66B0
    x"03",x"CC",x"01",x"40",x"DD",x"C7",x"CC",x"00", -- 0x66B8
    x"60",x"DD",x"C9",x"F6",x"FE",x"0B",x"8D",x"10", -- 0x66C0
    x"7E",x"E0",x"4D",x"50",x"A0",x"50",x"A0",x"26", -- 0x66C8
    x"05",x"F6",x"FE",x"0B",x"20",x"02",x"8D",x"36", -- 0x66D0
    x"0D",x"E6",x"27",x"13",x"8D",x"64",x"BD",x"E1", -- 0x66D8
    x"19",x"8E",x"20",x"00",x"E7",x"80",x"8C",x"A0", -- 0x66E0
    x"00",x"26",x"F9",x"BD",x"E0",x"FF",x"39",x"C6", -- 0x66E8
    x"4C",x"7E",x"AC",x"46",x"81",x"2C",x"10",x"21", -- 0x66F0
    x"19",x"06",x"27",x"09",x"8D",x"10",x"F7",x"FE", -- 0x66F8
    x"0A",x"9D",x"A5",x"27",x"08",x"BD",x"B2",x"6D", -- 0x6700
    x"8D",x"04",x"F7",x"FE",x"0B",x"39",x"BD",x"B7", -- 0x6708
    x"0B",x"C1",x"10",x"10",x"24",x"CD",x"33",x"39", -- 0x6710
    x"BD",x"E7",x"31",x"9D",x"A5",x"27",x"10",x"81", -- 0x6718
    x"29",x"27",x"0C",x"BD",x"B2",x"6D",x"81",x"2C", -- 0x6720
    x"27",x"05",x"BD",x"E7",x"0E",x"8D",x"0C",x"0E", -- 0x6728
    x"A5",x"F6",x"FE",x"0A",x"0D",x"C2",x"26",x"03", -- 0x6730
    x"F6",x"FE",x"0B",x"D7",x"B4",x"8D",x"03",x"D7", -- 0x6738
    x"B5",x"39",x"34",x"10",x"96",x"E6",x"80",x"01", -- 0x6740
    x"8E",x"E7",x"59",x"E4",x"86",x"96",x"E6",x"80", -- 0x6748
    x"01",x"8E",x"E7",x"5D",x"A6",x"86",x"3D",x"35", -- 0x6750
    x"90",x"03",x"0F",x"01",x"03",x"55",x"11",x"FF", -- 0x6758
    x"55",x"86",x"01",x"20",x"05",x"4F",x"10",x"21", -- 0x6760
    x"18",x"96",x"0D",x"E6",x"27",x"81",x"97",x"C2", -- 0x6768
    x"BD",x"B2",x"6A",x"BD",x"E7",x"AA",x"0D",x"C2", -- 0x6770
    x"26",x"05",x"BD",x"E7",x"31",x"20",x"03",x"BD", -- 0x6778
    x"E7",x"18",x"BD",x"B2",x"67",x"BD",x"E7",x"DA", -- 0x6780
    x"BD",x"E1",x"19",x"BD",x"E7",x"92",x"BD",x"E0", -- 0x6788
    x"FF",x"39",x"E6",x"84",x"34",x"04",x"1F",x"89", -- 0x6790
    x"43",x"A4",x"84",x"D4",x"B5",x"34",x"04",x"AA", -- 0x6798
    x"E0",x"A7",x"84",x"A0",x"E0",x"9A",x"DB",x"97", -- 0x67A0
    x"DB",x"39",x"BD",x"E7",x"B2",x"CE",x"00",x"BD", -- 0x67A8
    x"39",x"39",x"BD",x"B7",x"34",x"10",x"8E",x"00", -- 0x67B0
    x"BD",x"C1",x"C0",x"25",x"02",x"C6",x"BF",x"4F", -- 0x67B8
    x"ED",x"22",x"96",x"E6",x"81",x"02",x"2E",x"05", -- 0x67C0
    x"CC",x"01",x"3F",x"20",x"03",x"CC",x"02",x"7F", -- 0x67C8
    x"10",x"93",x"2B",x"25",x"02",x"DC",x"2B",x"ED", -- 0x67D0
    x"A4",x"39",x"8D",x"0A",x"6E",x"C4",x"E8",x"20", -- 0x67D8
    x"E8",x"3F",x"E7",x"FF",x"E8",x"20",x"CE",x"E7", -- 0x67E0
    x"DE",x"96",x"E6",x"80",x"01",x"48",x"EE",x"C6", -- 0x67E8
    x"39",x"80",x"40",x"20",x"10",x"08",x"04",x"02", -- 0x67F0
    x"01",x"C0",x"30",x"0C",x"03",x"F0",x"0F",x"34", -- 0x67F8
    x"44",x"D6",x"B9",x"96",x"C0",x"3D",x"C3",x"20", -- 0x6800
    x"00",x"1F",x"01",x"DC",x"BD",x"44",x"56",x"44", -- 0x6808
    x"56",x"44",x"56",x"30",x"8B",x"96",x"BE",x"84", -- 0x6810
    x"07",x"CE",x"E7",x"F1",x"A6",x"C6",x"35",x"C4", -- 0x6818
    x"34",x"44",x"D6",x"B9",x"96",x"C0",x"3D",x"C3", -- 0x6820
    x"20",x"00",x"1F",x"01",x"DC",x"BD",x"44",x"56", -- 0x6828
    x"44",x"56",x"30",x"8B",x"96",x"BE",x"84",x"03", -- 0x6830
    x"CE",x"E7",x"F9",x"A6",x"C6",x"35",x"C4",x"34", -- 0x6838
    x"44",x"D6",x"B9",x"96",x"C0",x"3D",x"C3",x"20", -- 0x6840
    x"00",x"1F",x"01",x"DC",x"BD",x"44",x"56",x"30", -- 0x6848
    x"8B",x"96",x"BE",x"84",x"01",x"CE",x"E7",x"FD", -- 0x6850
    x"A6",x"C6",x"35",x"C4",x"0D",x"E6",x"10",x"27", -- 0x6858
    x"FE",x"8D",x"BD",x"B2",x"6A",x"BD",x"E7",x"AA", -- 0x6860
    x"BD",x"B2",x"67",x"BD",x"E1",x"19",x"BD",x"E7", -- 0x6868
    x"DA",x"1F",x"89",x"E4",x"84",x"44",x"25",x"03", -- 0x6870
    x"54",x"20",x"FA",x"BD",x"B4",x"F3",x"BD",x"E0", -- 0x6878
    x"FF",x"39",x"0D",x"E6",x"10",x"27",x"FE",x"67", -- 0x6880
    x"10",x"21",x"17",x"74",x"81",x"28",x"27",x"09", -- 0x6888
    x"81",x"AC",x"27",x"05",x"C6",x"40",x"BD",x"B2", -- 0x6890
    x"6F",x"BD",x"E9",x"E1",x"9E",x"C3",x"9F",x"C7", -- 0x6898
    x"9E",x"C5",x"9F",x"C9",x"BD",x"B2",x"6D",x"81", -- 0x68A0
    x"BE",x"27",x"09",x"81",x"BD",x"10",x"26",x"C9", -- 0x68A8
    x"C6",x"C6",x"01",x"86",x"5F",x"34",x"04",x"9D", -- 0x68B0
    x"9F",x"BD",x"EA",x"0D",x"35",x"04",x"D7",x"C2", -- 0x68B8
    x"BD",x"E7",x"31",x"9D",x"A5",x"10",x"27",x"00", -- 0x68C0
    x"85",x"BD",x"B2",x"6D",x"C6",x"42",x"BD",x"B2", -- 0x68C8
    x"6F",x"26",x"18",x"8D",x"31",x"8D",x"5A",x"9E", -- 0x68D0
    x"BD",x"34",x"10",x"9E",x"C3",x"9F",x"BD",x"8D", -- 0x68D8
    x"50",x"35",x"10",x"9F",x"BD",x"9E",x"C5",x"9F", -- 0x68E0
    x"BF",x"20",x"1B",x"C6",x"46",x"BD",x"B2",x"6F", -- 0x68E8
    x"20",x"04",x"30",x"1F",x"9F",x"BF",x"BD",x"E9", -- 0x68F0
    x"06",x"9E",x"BF",x"9C",x"C5",x"27",x"06",x"24", -- 0x68F8
    x"F1",x"30",x"01",x"20",x"EF",x"39",x"9E",x"BD", -- 0x6900
    x"34",x"10",x"BD",x"E9",x"DB",x"24",x"04",x"9E", -- 0x6908
    x"C3",x"9F",x"BD",x"1F",x"02",x"31",x"21",x"BD", -- 0x6910
    x"E7",x"DA",x"35",x"40",x"DF",x"BD",x"17",x"00", -- 0x6918
    x"F5",x"97",x"D7",x"BD",x"E7",x"88",x"96",x"D7", -- 0x6920
    x"AD",x"C4",x"31",x"3F",x"26",x"F3",x"39",x"35", -- 0x6928
    x"06",x"DC",x"BF",x"34",x"06",x"BD",x"E9",x"CD", -- 0x6930
    x"24",x"04",x"9E",x"C5",x"9F",x"BF",x"1F",x"02", -- 0x6938
    x"31",x"21",x"BD",x"E7",x"DA",x"35",x"40",x"DF", -- 0x6940
    x"BF",x"17",x"00",x"D5",x"20",x"D3",x"10",x"8E", -- 0x6948
    x"E9",x"B8",x"BD",x"E9",x"CD",x"27",x"AF",x"24", -- 0x6950
    x"04",x"10",x"8E",x"E9",x"C6",x"34",x"06",x"CE", -- 0x6958
    x"E9",x"B1",x"BD",x"E9",x"DB",x"27",x"C8",x"24", -- 0x6960
    x"03",x"CE",x"E9",x"BF",x"10",x"A3",x"E4",x"35", -- 0x6968
    x"10",x"24",x"04",x"1E",x"32",x"1E",x"01",x"34", -- 0x6970
    x"46",x"34",x"06",x"44",x"56",x"25",x"09",x"11", -- 0x6978
    x"83",x"E9",x"B9",x"25",x"03",x"83",x"00",x"01", -- 0x6980
    x"34",x"16",x"BD",x"E7",x"E6",x"AD",x"C4",x"BD", -- 0x6988
    x"E7",x"88",x"AE",x"66",x"27",x"17",x"30",x"1F", -- 0x6990
    x"AF",x"66",x"AD",x"F8",x"08",x"EC",x"E4",x"E3", -- 0x6998
    x"62",x"ED",x"E4",x"A3",x"64",x"25",x"E6",x"ED", -- 0x69A0
    x"E4",x"AD",x"A4",x"20",x"E0",x"35",x"10",x"35", -- 0x69A8
    x"F6",x"9E",x"BD",x"30",x"01",x"9F",x"BD",x"39", -- 0x69B0
    x"9E",x"BF",x"30",x"01",x"9F",x"BF",x"39",x"9E", -- 0x69B8
    x"BD",x"30",x"1F",x"9F",x"BD",x"39",x"9E",x"BF", -- 0x69C0
    x"30",x"1F",x"9F",x"BF",x"39",x"DC",x"C5",x"93", -- 0x69C8
    x"BF",x"24",x"F9",x"34",x"01",x"40",x"50",x"82", -- 0x69D0
    x"00",x"35",x"81",x"DC",x"C3",x"93",x"BD",x"20", -- 0x69D8
    x"F0",x"9E",x"C7",x"9F",x"BD",x"9E",x"C9",x"9F", -- 0x69E0
    x"BF",x"81",x"AC",x"27",x"03",x"BD",x"EA",x"04", -- 0x69E8
    x"C6",x"AC",x"BD",x"B2",x"6F",x"BD",x"B2",x"6A", -- 0x69F0
    x"BD",x"B7",x"34",x"10",x"8E",x"00",x"C3",x"BD", -- 0x69F8
    x"E7",x"B9",x"20",x"06",x"BD",x"B2",x"6A",x"BD", -- 0x6A00
    x"E7",x"B2",x"7E",x"B2",x"67",x"BD",x"E7",x"AD", -- 0x6A08
    x"CE",x"00",x"C3",x"7E",x"E7",x"B0",x"CE",x"EA", -- 0x6A10
    x"25",x"D6",x"E6",x"C0",x"01",x"58",x"EE",x"C5", -- 0x6A18
    x"39",x"CE",x"EA",x"45",x"39",x"EA",x"34",x"EA", -- 0x6A20
    x"3D",x"EA",x"2D",x"EA",x"34",x"44",x"24",x"03", -- 0x6A28
    x"46",x"30",x"01",x"39",x"44",x"44",x"24",x"FB", -- 0x6A30
    x"86",x"C0",x"30",x"01",x"39",x"43",x"81",x"F0", -- 0x6A38
    x"26",x"02",x"30",x"01",x"39",x"D6",x"B9",x"3A", -- 0x6A40
    x"39",x"0D",x"E6",x"10",x"27",x"FC",x"A0",x"10", -- 0x6A48
    x"21",x"15",x"AD",x"81",x"40",x"26",x"02",x"9D", -- 0x6A50
    x"9F",x"BD",x"EB",x"60",x"BD",x"EA",x"04",x"BD", -- 0x6A58
    x"E7",x"AD",x"AE",x"C4",x"9F",x"CB",x"AE",x"42", -- 0x6A60
    x"9F",x"CD",x"BD",x"B2",x"6D",x"BD",x"B7",x"3D", -- 0x6A68
    x"CE",x"00",x"CF",x"AF",x"C4",x"BD",x"E7",x"B0", -- 0x6A70
    x"86",x"01",x"97",x"C2",x"BD",x"E7",x"18",x"8E", -- 0x6A78
    x"01",x"00",x"9D",x"A5",x"27",x"0F",x"BD",x"B2", -- 0x6A80
    x"6D",x"BD",x"B1",x"41",x"96",x"4F",x"8B",x"08", -- 0x6A88
    x"97",x"4F",x"BD",x"B7",x"40",x"96",x"E6",x"81", -- 0x6A90
    x"02",x"22",x"04",x"1F",x"10",x"30",x"8B",x"9F", -- 0x6A98
    x"D1",x"C6",x"01",x"D7",x"C2",x"D7",x"D8",x"BD", -- 0x6AA0
    x"EB",x"7B",x"34",x"06",x"BD",x"EB",x"7B",x"DD", -- 0x6AA8
    x"D9",x"35",x"06",x"34",x"06",x"9E",x"C3",x"9F", -- 0x6AB0
    x"BD",x"9E",x"C5",x"9F",x"BF",x"CE",x"EB",x"9B", -- 0x6AB8
    x"84",x"01",x"27",x"03",x"50",x"CB",x"08",x"58", -- 0x6AC0
    x"58",x"33",x"C5",x"34",x"40",x"BD",x"EB",x"BD", -- 0x6AC8
    x"35",x"40",x"33",x"5E",x"34",x"10",x"BD",x"EB", -- 0x6AD0
    x"BD",x"35",x"20",x"A6",x"E4",x"84",x"03",x"27", -- 0x6AD8
    x"06",x"81",x"03",x"27",x"02",x"1E",x"12",x"9F", -- 0x6AE0
    x"C3",x"1F",x"20",x"44",x"56",x"9E",x"D1",x"BD", -- 0x6AE8
    x"EB",x"CB",x"1F",x"20",x"4D",x"10",x"26",x"C9", -- 0x6AF0
    x"51",x"D7",x"C5",x"1F",x"30",x"97",x"C6",x"A6", -- 0x6AF8
    x"E4",x"81",x"02",x"25",x"0E",x"81",x"06",x"24", -- 0x6B00
    x"0A",x"DC",x"CB",x"93",x"C3",x"24",x"11",x"4F", -- 0x6B08
    x"5F",x"20",x"0D",x"DC",x"CB",x"D3",x"C3",x"25", -- 0x6B10
    x"05",x"10",x"93",x"D3",x"25",x"02",x"DC",x"D3", -- 0x6B18
    x"DD",x"C3",x"A6",x"E4",x"81",x"04",x"25",x"0A", -- 0x6B20
    x"DC",x"CD",x"93",x"C5",x"24",x"11",x"4F",x"5F", -- 0x6B28
    x"20",x"0D",x"DC",x"CD",x"D3",x"C5",x"25",x"05", -- 0x6B30
    x"10",x"93",x"D5",x"25",x"02",x"DC",x"D5",x"DD", -- 0x6B38
    x"C5",x"0D",x"D8",x"26",x"03",x"17",x"FE",x"06", -- 0x6B40
    x"35",x"06",x"04",x"D8",x"25",x"05",x"10",x"93", -- 0x6B48
    x"D9",x"27",x"0C",x"5C",x"C1",x"08",x"26",x"04", -- 0x6B50
    x"4C",x"5F",x"84",x"07",x"7E",x"EA",x"B3",x"39", -- 0x6B58
    x"CE",x"00",x"D3",x"8E",x"02",x"7F",x"AF",x"C4", -- 0x6B60
    x"96",x"E6",x"81",x"02",x"2E",x"05",x"8E",x"01", -- 0x6B68
    x"3F",x"AF",x"C4",x"8E",x"00",x"BF",x"AF",x"42", -- 0x6B70
    x"7E",x"E7",x"B0",x"5F",x"9D",x"A5",x"27",x"11", -- 0x6B78
    x"BD",x"B2",x"6D",x"BD",x"B1",x"41",x"96",x"4F", -- 0x6B80
    x"8B",x"06",x"97",x"4F",x"BD",x"B7",x"0E",x"C4", -- 0x6B88
    x"3F",x"1F",x"98",x"C4",x"07",x"44",x"44",x"44", -- 0x6B90
    x"39",x"00",x"00",x"00",x"01",x"FE",x"C5",x"19", -- 0x6B98
    x"19",x"FB",x"16",x"31",x"F2",x"F4",x"FB",x"4A", -- 0x6BA0
    x"51",x"EC",x"84",x"61",x"F9",x"E1",x"C7",x"78", -- 0x6BA8
    x"AE",x"D4",x"DC",x"8E",x"3B",x"C5",x"E5",x"A2", -- 0x6BB0
    x"69",x"B5",x"06",x"B5",x"06",x"9E",x"CF",x"EC", -- 0x6BB8
    x"C4",x"27",x"07",x"83",x"00",x"01",x"8D",x"03", -- 0x6BC0
    x"1F",x"21",x"39",x"34",x"76",x"6F",x"64",x"A6", -- 0x6BC8
    x"63",x"3D",x"ED",x"66",x"EC",x"61",x"3D",x"EB", -- 0x6BD0
    x"66",x"89",x"00",x"ED",x"65",x"E6",x"E4",x"A6", -- 0x6BD8
    x"63",x"3D",x"E3",x"65",x"ED",x"65",x"24",x"02", -- 0x6BE0
    x"6C",x"64",x"A6",x"E4",x"E6",x"62",x"3D",x"E3", -- 0x6BE8
    x"64",x"ED",x"64",x"35",x"F6",x"0D",x"E6",x"10", -- 0x6BF0
    x"27",x"FA",x"F4",x"10",x"21",x"14",x"01",x"81", -- 0x6BF8
    x"40",x"26",x"02",x"9D",x"9F",x"BD",x"EA",x"04", -- 0x6C00
    x"BD",x"E7",x"AD",x"86",x"01",x"97",x"C2",x"BD", -- 0x6C08
    x"E7",x"18",x"DC",x"B4",x"34",x"06",x"9D",x"A5", -- 0x6C10
    x"27",x"03",x"BD",x"E7",x"18",x"96",x"B5",x"97", -- 0x6C18
    x"D8",x"35",x"06",x"DD",x"B4",x"BD",x"E1",x"19", -- 0x6C20
    x"4F",x"34",x"56",x"BD",x"EB",x"60",x"BD",x"E7", -- 0x6C28
    x"E6",x"DF",x"D9",x"BD",x"EC",x"BE",x"27",x"0F", -- 0x6C30
    x"BD",x"ED",x"01",x"86",x"01",x"97",x"D7",x"BD", -- 0x6C38
    x"ED",x"2E",x"00",x"D7",x"BD",x"ED",x"2E",x"10", -- 0x6C40
    x"DF",x"DC",x"0D",x"DB",x"26",x"03",x"10",x"DE", -- 0x6C48
    x"DC",x"35",x"56",x"0F",x"DB",x"10",x"DF",x"DC", -- 0x6C50
    x"30",x"01",x"9F",x"BD",x"DF",x"D1",x"97",x"D7", -- 0x6C58
    x"27",x"58",x"2B",x"06",x"5C",x"D1",x"D6",x"23", -- 0x6C60
    x"05",x"5F",x"5D",x"27",x"DD",x"5A",x"D7",x"C0", -- 0x6C68
    x"BD",x"EC",x"BE",x"27",x"11",x"10",x"83",x"00", -- 0x6C70
    x"03",x"25",x"05",x"30",x"1E",x"BD",x"ED",x"15", -- 0x6C78
    x"BD",x"ED",x"01",x"BD",x"ED",x"2E",x"43",x"53", -- 0x6C80
    x"D3",x"D1",x"DD",x"D1",x"2F",x"17",x"BD",x"E9", -- 0x6C88
    x"B1",x"BD",x"EC",x"F1",x"26",x"05",x"CC",x"FF", -- 0x6C90
    x"FF",x"20",x"ED",x"BD",x"E9",x"BF",x"BD",x"ED", -- 0x6C98
    x"3A",x"8D",x"24",x"20",x"DE",x"BD",x"E9",x"B1", -- 0x6CA0
    x"30",x"8B",x"9F",x"BD",x"43",x"53",x"83",x"00", -- 0x6CA8
    x"01",x"2F",x"04",x"1F",x"01",x"8D",x"5E",x"7E", -- 0x6CB0
    x"EC",x"4A",x"BD",x"E0",x"FF",x"39",x"BD",x"ED", -- 0x6CB8
    x"3A",x"10",x"8E",x"E9",x"BF",x"20",x"06",x"10", -- 0x6CC0
    x"8E",x"E9",x"B1",x"AD",x"A4",x"DE",x"8A",x"9E", -- 0x6CC8
    x"BD",x"2B",x"17",x"9C",x"D3",x"22",x"13",x"34", -- 0x6CD0
    x"60",x"8D",x"16",x"27",x"0B",x"BD",x"E7",x"92", -- 0x6CD8
    x"35",x"60",x"33",x"41",x"AD",x"A4",x"20",x"E9", -- 0x6CE0
    x"35",x"60",x"1F",x"30",x"1F",x"01",x"93",x"8A", -- 0x6CE8
    x"39",x"AD",x"9F",x"00",x"D9",x"1F",x"89",x"D4", -- 0x6CF0
    x"D8",x"34",x"06",x"A4",x"84",x"A1",x"61",x"35", -- 0x6CF8
    x"86",x"DD",x"CD",x"10",x"9E",x"C3",x"8D",x"32", -- 0x6D00
    x"10",x"9F",x"BD",x"8D",x"BA",x"9E",x"CD",x"30", -- 0x6D08
    x"8B",x"C3",x"00",x"01",x"39",x"DD",x"CB",x"35", -- 0x6D10
    x"20",x"DC",x"BD",x"34",x"16",x"96",x"D7",x"40", -- 0x6D18
    x"D6",x"C0",x"34",x"06",x"34",x"20",x"C6",x"06", -- 0x6D20
    x"BD",x"ED",x"3F",x"DC",x"CB",x"39",x"DD",x"CB", -- 0x6D28
    x"35",x"20",x"DC",x"C3",x"34",x"16",x"96",x"D7", -- 0x6D30
    x"20",x"E6",x"9E",x"BD",x"9F",x"C3",x"39",x"50", -- 0x6D38
    x"32",x"E5",x"11",x"8C",x"BF",x"F1",x"10",x"25", -- 0x6D40
    x"00",x"04",x"50",x"32",x"E5",x"39",x"10",x"CE", -- 0x6D48
    x"DF",x"FD",x"BD",x"E0",x"FF",x"7E",x"AC",x"44", -- 0x6D50
    x"BD",x"B7",x"3D",x"10",x"21",x"12",x"A1",x"8C", -- 0x6D58
    x"00",x"FF",x"10",x"22",x"C6",x"E4",x"9F",x"D1", -- 0x6D60
    x"27",x"08",x"BD",x"B2",x"6D",x"BD",x"B7",x"3D", -- 0x6D68
    x"9F",x"D3",x"BD",x"E0",x"CB",x"BD",x"E1",x"19", -- 0x6D70
    x"DC",x"D1",x"5D",x"26",x"08",x"CC",x"FF",x"FF", -- 0x6D78
    x"FD",x"C0",x"00",x"20",x"38",x"10",x"8E",x"C0", -- 0x6D80
    x"00",x"EC",x"A4",x"10",x"83",x"FF",x"FF",x"26", -- 0x6D88
    x"04",x"8D",x"31",x"20",x"1B",x"D6",x"D2",x"E1", -- 0x6D90
    x"22",x"27",x"37",x"EE",x"A4",x"27",x"04",x"1F", -- 0x6D98
    x"32",x"20",x"F4",x"1F",x"23",x"EC",x"23",x"31", -- 0x6DA0
    x"25",x"31",x"AB",x"8D",x"17",x"10",x"AF",x"C4", -- 0x6DA8
    x"CC",x"00",x"00",x"ED",x"A4",x"D6",x"D2",x"E7", -- 0x6DB0
    x"22",x"DC",x"D3",x"ED",x"23",x"BD",x"E0",x"FF", -- 0x6DB8
    x"BD",x"E0",x"97",x"39",x"1F",x"21",x"30",x"05", -- 0x6DC0
    x"DC",x"D3",x"30",x"8B",x"8C",x"DF",x"00",x"22", -- 0x6DC8
    x"05",x"39",x"C6",x"12",x"20",x"02",x"C6",x"0C", -- 0x6DD0
    x"10",x"CE",x"DF",x"FD",x"BD",x"E0",x"FF",x"BD", -- 0x6DD8
    x"E0",x"97",x"7E",x"AC",x"46",x"8E",x"EE",x"C0", -- 0x6DE0
    x"9F",x"D5",x"5F",x"20",x"07",x"8E",x"EE",x"EF", -- 0x6DE8
    x"9F",x"D5",x"C6",x"01",x"0D",x"E6",x"10",x"27", -- 0x6DF0
    x"F8",x"F5",x"10",x"21",x"12",x"02",x"D7",x"D8", -- 0x6DF8
    x"81",x"40",x"26",x"02",x"9D",x"9F",x"BD",x"E9", -- 0x6E00
    x"E1",x"BD",x"B2",x"6D",x"BD",x"B7",x"0B",x"D7", -- 0x6E08
    x"D3",x"0F",x"D4",x"9D",x"A5",x"27",x"21",x"03", -- 0x6E10
    x"D4",x"BD",x"B2",x"6D",x"0D",x"D8",x"26",x"03", -- 0x6E18
    x"16",x"C4",x"54",x"C6",x"05",x"8E",x"EE",x"E0", -- 0x6E20
    x"EE",x"81",x"A1",x"80",x"27",x"06",x"5A",x"26", -- 0x6E28
    x"F7",x"7E",x"B2",x"77",x"DF",x"D5",x"9D",x"9F", -- 0x6E30
    x"BD",x"E0",x"CB",x"BD",x"E1",x"19",x"D6",x"D3", -- 0x6E38
    x"BD",x"EF",x"18",x"DC",x"BD",x"10",x"93",x"C3", -- 0x6E40
    x"2F",x"06",x"9E",x"C3",x"9F",x"BD",x"DD",x"C3", -- 0x6E48
    x"DC",x"BF",x"10",x"93",x"C5",x"2F",x"06",x"9E", -- 0x6E50
    x"C5",x"9F",x"BF",x"DD",x"C5",x"96",x"E6",x"C6", -- 0x6E58
    x"F8",x"81",x"03",x"27",x"08",x"C6",x"FC",x"81", -- 0x6E60
    x"02",x"26",x"02",x"C6",x"FE",x"1F",x"98",x"94", -- 0x6E68
    x"BE",x"97",x"BE",x"D4",x"C4",x"D7",x"C4",x"BD", -- 0x6E70
    x"E9",x"DB",x"DD",x"C3",x"BD",x"E9",x"CD",x"C3", -- 0x6E78
    x"00",x"01",x"DD",x"C5",x"96",x"E6",x"81",x"02", -- 0x6E80
    x"27",x"0C",x"81",x"03",x"26",x"04",x"04",x"C3", -- 0x6E88
    x"06",x"C4",x"04",x"C3",x"06",x"C4",x"04",x"C3", -- 0x6E90
    x"06",x"C4",x"DC",x"C3",x"C3",x"00",x"01",x"DD", -- 0x6E98
    x"C3",x"BD",x"E7",x"DA",x"10",x"9E",x"D5",x"D6", -- 0x6EA0
    x"C4",x"34",x"10",x"AD",x"A4",x"5A",x"26",x"FB", -- 0x6EA8
    x"35",x"10",x"BD",x"EA",x"45",x"0A",x"C6",x"26", -- 0x6EB0
    x"EE",x"BD",x"E0",x"FF",x"BD",x"E0",x"97",x"39", -- 0x6EB8
    x"A6",x"80",x"8D",x"03",x"A7",x"C4",x"39",x"DE", -- 0x6EC0
    x"CF",x"33",x"41",x"DF",x"CF",x"11",x"93",x"D1", -- 0x6EC8
    x"22",x"01",x"39",x"10",x"CE",x"DF",x"FD",x"BD", -- 0x6ED0
    x"E0",x"FF",x"BD",x"E0",x"97",x"7E",x"B4",x"4A", -- 0x6ED8
    x"EE",x"EF",x"BD",x"EE",x"F6",x"BE",x"EF",x"07", -- 0x6EE0
    x"B1",x"EE",x"FE",x"B0",x"EF",x"10",x"A8",x"8D", -- 0x6EE8
    x"D6",x"A6",x"C4",x"A7",x"80",x"39",x"8D",x"CF", -- 0x6EF0
    x"A6",x"C4",x"43",x"A7",x"80",x"39",x"8D",x"C7", -- 0x6EF8
    x"A6",x"C4",x"A4",x"84",x"A7",x"80",x"39",x"8D", -- 0x6F00
    x"BE",x"A6",x"C4",x"AA",x"84",x"A7",x"80",x"39", -- 0x6F08
    x"8D",x"B5",x"A6",x"84",x"43",x"A7",x"80",x"39", -- 0x6F10
    x"10",x"8E",x"C0",x"00",x"A6",x"A4",x"81",x"FF", -- 0x6F18
    x"26",x"0A",x"7E",x"EE",x"D3",x"10",x"AE",x"A4", -- 0x6F20
    x"10",x"27",x"FF",x"A7",x"E1",x"22",x"26",x"F5", -- 0x6F28
    x"EC",x"23",x"31",x"24",x"10",x"9F",x"CF",x"31", -- 0x6F30
    x"21",x"31",x"AB",x"10",x"9F",x"D1",x"39",x"0D", -- 0x6F38
    x"E6",x"10",x"27",x"F7",x"AA",x"10",x"21",x"10", -- 0x6F40
    x"B7",x"BD",x"B2",x"6A",x"BD",x"E7",x"B2",x"BD", -- 0x6F48
    x"B2",x"67",x"BD",x"B2",x"6D",x"BD",x"B1",x"56", -- 0x6F50
    x"0D",x"06",x"26",x"06",x"BD",x"BD",x"D9",x"BD", -- 0x6F58
    x"B5",x"16",x"BD",x"B6",x"57",x"F7",x"FE",x"18", -- 0x6F60
    x"10",x"8E",x"FE",x"19",x"5A",x"2B",x"06",x"A6", -- 0x6F68
    x"80",x"A7",x"A0",x"20",x"F7",x"96",x"E6",x"C6", -- 0x6F70
    x"28",x"81",x"03",x"25",x"02",x"C6",x"50",x"4F", -- 0x6F78
    x"93",x"BD",x"2B",x"7D",x"F1",x"FE",x"18",x"22", -- 0x6F80
    x"05",x"F7",x"FE",x"18",x"27",x"73",x"86",x"17", -- 0x6F88
    x"91",x"C0",x"2C",x"02",x"97",x"C0",x"BD",x"F0", -- 0x6F90
    x"8C",x"BD",x"E7",x"DA",x"10",x"8E",x"FE",x"19", -- 0x6F98
    x"F6",x"FE",x"18",x"A6",x"A4",x"84",x"7F",x"80", -- 0x6FA0
    x"20",x"2A",x"02",x"86",x"00",x"A7",x"A0",x"5A", -- 0x6FA8
    x"2E",x"F1",x"96",x"E6",x"4A",x"48",x"10",x"8E", -- 0x6FB0
    x"F0",x"02",x"10",x"AE",x"A6",x"10",x"9F",x"D1", -- 0x6FB8
    x"86",x"08",x"97",x"D3",x"10",x"8E",x"FE",x"19", -- 0x6FC0
    x"CE",x"F0",x"9D",x"F6",x"FE",x"0A",x"BD",x"E7", -- 0x6FC8
    x"42",x"D7",x"B5",x"BD",x"E1",x"19",x"B6",x"FE", -- 0x6FD0
    x"18",x"34",x"32",x"E6",x"A0",x"4F",x"58",x"58", -- 0x6FD8
    x"49",x"58",x"49",x"A6",x"CB",x"AD",x"9F",x"00", -- 0x6FE0
    x"D1",x"7A",x"FE",x"18",x"2E",x"ED",x"35",x"32", -- 0x6FE8
    x"0A",x"D3",x"27",x"0A",x"B7",x"FE",x"18",x"33", -- 0x6FF0
    x"41",x"BD",x"EA",x"45",x"20",x"DB",x"BD",x"E0", -- 0x6FF8
    x"FF",x"39",x"F0",x"1A",x"F0",x"45",x"F0",x"0A", -- 0x7000
    x"F0",x"1A",x"34",x"02",x"43",x"A4",x"84",x"A7", -- 0x7008
    x"84",x"35",x"02",x"94",x"B5",x"AA",x"84",x"A7", -- 0x7010
    x"80",x"39",x"34",x"20",x"10",x"8E",x"F0",x"35", -- 0x7018
    x"1F",x"89",x"44",x"44",x"44",x"44",x"A6",x"A6", -- 0x7020
    x"BD",x"F0",x"0A",x"C4",x"0F",x"A6",x"A5",x"BD", -- 0x7028
    x"F0",x"0A",x"35",x"20",x"39",x"00",x"03",x"0C", -- 0x7030
    x"0F",x"30",x"33",x"3C",x"3F",x"C0",x"C3",x"CC", -- 0x7038
    x"CF",x"F0",x"F3",x"FC",x"FF",x"34",x"22",x"10", -- 0x7040
    x"8E",x"F0",x"6C",x"44",x"44",x"44",x"44",x"48", -- 0x7048
    x"EC",x"A6",x"BD",x"F0",x"0A",x"1F",x"98",x"BD", -- 0x7050
    x"F0",x"0A",x"35",x"02",x"84",x"0F",x"48",x"EC", -- 0x7058
    x"A6",x"BD",x"F0",x"0A",x"1F",x"98",x"BD",x"F0", -- 0x7060
    x"0A",x"35",x"20",x"39",x"00",x"00",x"00",x"0F", -- 0x7068
    x"00",x"F0",x"00",x"FF",x"0F",x"00",x"0F",x"0F", -- 0x7070
    x"0F",x"F0",x"0F",x"FF",x"F0",x"00",x"F0",x"0F", -- 0x7078
    x"F0",x"F0",x"F0",x"FF",x"FF",x"00",x"FF",x"0F", -- 0x7080
    x"FF",x"F0",x"FF",x"FF",x"DC",x"BD",x"58",x"58", -- 0x7088
    x"49",x"58",x"49",x"DD",x"BD",x"96",x"C0",x"48", -- 0x7090
    x"48",x"48",x"97",x"C0",x"39",x"00",x"00",x"00", -- 0x7098
    x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10", -- 0x70A0
    x"10",x"10",x"00",x"10",x"00",x"28",x"28",x"28", -- 0x70A8
    x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"7C", -- 0x70B0
    x"28",x"7C",x"28",x"28",x"00",x"10",x"3C",x"50", -- 0x70B8
    x"38",x"14",x"78",x"10",x"00",x"60",x"64",x"08", -- 0x70C0
    x"10",x"20",x"4C",x"0C",x"00",x"20",x"50",x"50", -- 0x70C8
    x"20",x"54",x"48",x"34",x"00",x"10",x"10",x"20", -- 0x70D0
    x"00",x"00",x"00",x"00",x"00",x"08",x"10",x"20", -- 0x70D8
    x"20",x"20",x"10",x"08",x"00",x"20",x"10",x"08", -- 0x70E0
    x"08",x"08",x"10",x"20",x"00",x"00",x"10",x"54", -- 0x70E8
    x"38",x"38",x"54",x"10",x"00",x"00",x"10",x"10", -- 0x70F0
    x"7C",x"10",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x70F8
    x"00",x"00",x"10",x"10",x"20",x"00",x"00",x"00", -- 0x7100
    x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7108
    x"00",x"00",x"00",x"10",x"00",x"00",x"04",x"08", -- 0x7110
    x"10",x"20",x"40",x"00",x"00",x"38",x"44",x"4C", -- 0x7118
    x"54",x"64",x"44",x"38",x"00",x"10",x"30",x"10", -- 0x7120
    x"10",x"10",x"10",x"38",x"00",x"38",x"44",x"04", -- 0x7128
    x"38",x"40",x"40",x"7C",x"00",x"38",x"44",x"04", -- 0x7130
    x"08",x"04",x"44",x"38",x"00",x"08",x"18",x"28", -- 0x7138
    x"48",x"7C",x"08",x"08",x"00",x"7C",x"40",x"78", -- 0x7140
    x"04",x"04",x"44",x"38",x"00",x"38",x"40",x"40", -- 0x7148
    x"78",x"44",x"44",x"38",x"00",x"7C",x"04",x"08", -- 0x7150
    x"10",x"20",x"40",x"40",x"00",x"38",x"44",x"44", -- 0x7158
    x"38",x"44",x"44",x"38",x"00",x"38",x"44",x"44", -- 0x7160
    x"38",x"04",x"04",x"38",x"00",x"00",x"00",x"10", -- 0x7168
    x"00",x"00",x"10",x"00",x"00",x"00",x"00",x"10", -- 0x7170
    x"00",x"00",x"10",x"10",x"20",x"08",x"10",x"20", -- 0x7178
    x"40",x"20",x"10",x"08",x"00",x"00",x"00",x"7C", -- 0x7180
    x"00",x"7C",x"00",x"00",x"00",x"20",x"10",x"08", -- 0x7188
    x"04",x"08",x"10",x"20",x"00",x"38",x"44",x"04", -- 0x7190
    x"08",x"10",x"00",x"10",x"00",x"38",x"44",x"04", -- 0x7198
    x"34",x"4C",x"4C",x"38",x"00",x"10",x"28",x"44", -- 0x71A0
    x"44",x"7C",x"44",x"44",x"00",x"78",x"24",x"24", -- 0x71A8
    x"38",x"24",x"24",x"78",x"00",x"38",x"44",x"40", -- 0x71B0
    x"40",x"40",x"44",x"38",x"00",x"78",x"24",x"24", -- 0x71B8
    x"24",x"24",x"24",x"78",x"00",x"7C",x"40",x"40", -- 0x71C0
    x"70",x"40",x"40",x"7C",x"00",x"7C",x"40",x"40", -- 0x71C8
    x"70",x"40",x"40",x"40",x"00",x"38",x"44",x"40", -- 0x71D0
    x"40",x"4C",x"44",x"38",x"00",x"44",x"44",x"44", -- 0x71D8
    x"7C",x"44",x"44",x"44",x"00",x"38",x"10",x"10", -- 0x71E0
    x"10",x"10",x"10",x"38",x"00",x"04",x"04",x"04", -- 0x71E8
    x"04",x"04",x"44",x"38",x"00",x"44",x"48",x"50", -- 0x71F0
    x"60",x"50",x"48",x"44",x"00",x"40",x"40",x"40", -- 0x71F8
    x"40",x"40",x"40",x"7C",x"00",x"44",x"6C",x"54", -- 0x7200
    x"54",x"44",x"44",x"44",x"00",x"44",x"44",x"64", -- 0x7208
    x"54",x"4C",x"44",x"44",x"00",x"38",x"44",x"44", -- 0x7210
    x"44",x"44",x"44",x"38",x"00",x"78",x"44",x"44", -- 0x7218
    x"78",x"40",x"40",x"40",x"00",x"38",x"44",x"44", -- 0x7220
    x"44",x"54",x"48",x"34",x"00",x"78",x"44",x"44", -- 0x7228
    x"78",x"50",x"48",x"44",x"00",x"38",x"44",x"40", -- 0x7230
    x"38",x"04",x"44",x"38",x"00",x"7C",x"10",x"10", -- 0x7238
    x"10",x"10",x"10",x"10",x"00",x"44",x"44",x"44", -- 0x7240
    x"44",x"44",x"44",x"38",x"00",x"44",x"44",x"44", -- 0x7248
    x"28",x"28",x"10",x"10",x"00",x"44",x"44",x"44", -- 0x7250
    x"44",x"54",x"6C",x"44",x"00",x"44",x"44",x"28", -- 0x7258
    x"10",x"28",x"44",x"44",x"00",x"44",x"44",x"28", -- 0x7260
    x"10",x"10",x"10",x"10",x"00",x"7C",x"04",x"08", -- 0x7268
    x"10",x"20",x"40",x"7C",x"00",x"38",x"20",x"20", -- 0x7270
    x"20",x"20",x"20",x"38",x"00",x"00",x"40",x"20", -- 0x7278
    x"10",x"08",x"04",x"00",x"00",x"38",x"08",x"08", -- 0x7280
    x"08",x"08",x"08",x"38",x"00",x"10",x"38",x"54", -- 0x7288
    x"10",x"10",x"10",x"10",x"00",x"00",x"10",x"20", -- 0x7290
    x"7C",x"20",x"10",x"00",x"00",x"10",x"28",x"44", -- 0x7298
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38", -- 0x72A0
    x"04",x"3C",x"44",x"3C",x"00",x"40",x"40",x"58", -- 0x72A8
    x"64",x"44",x"64",x"58",x"00",x"00",x"00",x"38", -- 0x72B0
    x"44",x"40",x"44",x"38",x"00",x"04",x"04",x"34", -- 0x72B8
    x"4C",x"44",x"4C",x"34",x"00",x"00",x"00",x"38", -- 0x72C0
    x"44",x"7C",x"40",x"38",x"00",x"08",x"14",x"10", -- 0x72C8
    x"38",x"10",x"10",x"10",x"00",x"00",x"00",x"34", -- 0x72D0
    x"4C",x"4C",x"34",x"04",x"38",x"40",x"40",x"58", -- 0x72D8
    x"64",x"44",x"44",x"44",x"00",x"00",x"10",x"00", -- 0x72E0
    x"30",x"10",x"10",x"38",x"00",x"00",x"04",x"00", -- 0x72E8
    x"04",x"04",x"04",x"44",x"38",x"40",x"40",x"48", -- 0x72F0
    x"50",x"60",x"50",x"48",x"00",x"30",x"10",x"10", -- 0x72F8
    x"10",x"10",x"10",x"38",x"00",x"00",x"00",x"68", -- 0x7300
    x"54",x"54",x"54",x"54",x"00",x"00",x"00",x"58", -- 0x7308
    x"64",x"44",x"44",x"44",x"00",x"00",x"00",x"38", -- 0x7310
    x"44",x"44",x"44",x"38",x"00",x"00",x"00",x"78", -- 0x7318
    x"44",x"44",x"78",x"40",x"40",x"00",x"00",x"3C", -- 0x7320
    x"44",x"44",x"3C",x"04",x"04",x"00",x"00",x"58", -- 0x7328
    x"64",x"40",x"40",x"40",x"00",x"00",x"00",x"3C", -- 0x7330
    x"40",x"38",x"04",x"78",x"00",x"20",x"20",x"70", -- 0x7338
    x"20",x"20",x"24",x"18",x"00",x"00",x"00",x"44", -- 0x7340
    x"44",x"44",x"4C",x"34",x"00",x"00",x"00",x"44", -- 0x7348
    x"44",x"44",x"28",x"10",x"00",x"00",x"00",x"44", -- 0x7350
    x"54",x"54",x"28",x"28",x"00",x"00",x"00",x"44", -- 0x7358
    x"28",x"10",x"28",x"44",x"00",x"00",x"00",x"44", -- 0x7360
    x"44",x"44",x"3C",x"04",x"38",x"00",x"00",x"7C", -- 0x7368
    x"08",x"10",x"20",x"7C",x"00",x"08",x"10",x"10", -- 0x7370
    x"20",x"10",x"10",x"08",x"00",x"10",x"10",x"10", -- 0x7378
    x"00",x"10",x"10",x"10",x"00",x"20",x"10",x"10", -- 0x7380
    x"08",x"10",x"10",x"20",x"00",x"20",x"54",x"08", -- 0x7388
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7390
    x"00",x"00",x"00",x"7C",x"00",x"0D",x"E6",x"10", -- 0x7398
    x"27",x"F3",x"4C",x"10",x"21",x"0C",x"59",x"8E", -- 0x73A0
    x"00",x"00",x"C6",x"01",x"34",x"14",x"D7",x"C2", -- 0x73A8
    x"9F",x"D5",x"BD",x"E7",x"31",x"BD",x"B1",x"56", -- 0x73B0
    x"BD",x"B6",x"54",x"20",x"08",x"BD",x"F5",x"91", -- 0x73B8
    x"7E",x"F5",x"A7",x"35",x"14",x"D7",x"D8",x"27", -- 0x73C0
    x"FA",x"9F",x"D9",x"10",x"27",x"01",x"01",x"0D", -- 0x73C8
    x"D8",x"27",x"F0",x"BD",x"F5",x"91",x"81",x"3B", -- 0x73D0
    x"27",x"F5",x"81",x"27",x"27",x"F1",x"81",x"4E", -- 0x73D8
    x"26",x"04",x"03",x"D5",x"20",x"E9",x"81",x"42", -- 0x73E0
    x"26",x"04",x"03",x"D6",x"20",x"E1",x"81",x"58", -- 0x73E8
    x"10",x"27",x"00",x"AD",x"81",x"4D",x"10",x"27", -- 0x73F0
    x"01",x"52",x"34",x"02",x"C6",x"01",x"0F",x"D3", -- 0x73F8
    x"D7",x"D4",x"0D",x"D8",x"27",x"11",x"BD",x"F5", -- 0x7400
    x"91",x"BD",x"B3",x"A2",x"34",x"01",x"BD",x"F5", -- 0x7408
    x"F2",x"35",x"01",x"24",x"02",x"8D",x"A6",x"35", -- 0x7410
    x"02",x"81",x"43",x"27",x"28",x"81",x"41",x"27", -- 0x7418
    x"30",x"81",x"53",x"27",x"37",x"81",x"55",x"27", -- 0x7420
    x"6D",x"81",x"44",x"27",x"65",x"81",x"4C",x"27", -- 0x7428
    x"5B",x"81",x"52",x"27",x"50",x"80",x"45",x"27", -- 0x7430
    x"3A",x"4A",x"27",x"31",x"4A",x"27",x"3E",x"4A", -- 0x7438
    x"27",x"25",x"7E",x"B4",x"4A",x"BD",x"E7",x"11", -- 0x7440
    x"F7",x"FE",x"0A",x"BD",x"E7",x"31",x"16",x"FF", -- 0x7448
    x"7E",x"C1",x"04",x"10",x"24",x"BF",x"F3",x"D7", -- 0x7450
    x"E8",x"16",x"FF",x"73",x"C1",x"3F",x"10",x"24", -- 0x7458
    x"BF",x"E8",x"D7",x"E9",x"16",x"FF",x"68",x"96", -- 0x7460
    x"D3",x"8D",x"61",x"20",x"02",x"96",x"D3",x"1F", -- 0x7468
    x"01",x"20",x"61",x"96",x"D3",x"1F",x"01",x"8D", -- 0x7470
    x"53",x"1E",x"01",x"20",x"57",x"96",x"D3",x"1F", -- 0x7478
    x"01",x"8D",x"49",x"20",x"4F",x"96",x"D3",x"8E", -- 0x7480
    x"00",x"00",x"20",x"48",x"96",x"D3",x"8D",x"3C", -- 0x7488
    x"20",x"F5",x"96",x"D3",x"20",x"04",x"96",x"D3", -- 0x7490
    x"8D",x"32",x"8E",x"00",x"00",x"1E",x"10",x"20", -- 0x7498
    x"33",x"BD",x"F6",x"11",x"C6",x"02",x"BD",x"AC", -- 0x74A0
    x"33",x"D6",x"D8",x"9E",x"D9",x"34",x"14",x"7E", -- 0x74A8
    x"F3",x"B8",x"D6",x"E9",x"27",x"1B",x"4F",x"1E", -- 0x74B0
    x"01",x"A7",x"E2",x"2A",x"02",x"8D",x"0D",x"BD", -- 0x74B8
    x"EB",x"CB",x"1F",x"30",x"44",x"56",x"44",x"56", -- 0x74C0
    x"6D",x"E0",x"2A",x"04",x"40",x"50",x"82",x"00", -- 0x74C8
    x"39",x"1F",x"10",x"39",x"34",x"06",x"8D",x"DA", -- 0x74D0
    x"35",x"10",x"34",x"06",x"8D",x"D4",x"35",x"10", -- 0x74D8
    x"10",x"9E",x"E8",x"34",x"20",x"6D",x"E4",x"27", -- 0x74E0
    x"08",x"1E",x"10",x"8D",x"DF",x"6A",x"E4",x"20", -- 0x74E8
    x"F4",x"35",x"20",x"CE",x"00",x"00",x"D3",x"C7", -- 0x74F0
    x"2B",x"02",x"1F",x"03",x"1F",x"10",x"8E",x"00", -- 0x74F8
    x"00",x"D3",x"C9",x"2B",x"02",x"1F",x"01",x"11", -- 0x7500
    x"83",x"02",x"80",x"25",x"03",x"CE",x"02",x"7F", -- 0x7508
    x"96",x"E6",x"81",x"02",x"2E",x"09",x"11",x"83", -- 0x7510
    x"01",x"40",x"25",x"03",x"CE",x"01",x"3F",x"8C", -- 0x7518
    x"00",x"C0",x"25",x"03",x"8E",x"00",x"BF",x"DC", -- 0x7520
    x"C7",x"DD",x"BD",x"DC",x"C9",x"DD",x"BF",x"9F", -- 0x7528
    x"C5",x"DF",x"C3",x"0D",x"D5",x"26",x"04",x"9F", -- 0x7530
    x"C9",x"DF",x"C7",x"BD",x"EA",x"0D",x"0D",x"D6", -- 0x7538
    x"26",x"03",x"BD",x"E9",x"4E",x"0F",x"D5",x"0F", -- 0x7540
    x"D6",x"7E",x"F3",x"CF",x"BD",x"F5",x"91",x"34", -- 0x7548
    x"02",x"BD",x"F5",x"78",x"34",x"06",x"BD",x"F5", -- 0x7550
    x"91",x"81",x"2C",x"10",x"26",x"BE",x"EB",x"BD", -- 0x7558
    x"F5",x"75",x"1F",x"01",x"35",x"40",x"35",x"02", -- 0x7560
    x"81",x"2B",x"27",x"04",x"81",x"2D",x"26",x"97", -- 0x7568
    x"1F",x"30",x"7E",x"F4",x"D4",x"BD",x"F5",x"91", -- 0x7570
    x"81",x"2B",x"27",x"07",x"81",x"2D",x"27",x"04", -- 0x7578
    x"BD",x"F5",x"F2",x"4F",x"34",x"02",x"BD",x"F3", -- 0x7580
    x"BD",x"6D",x"E0",x"27",x"03",x"50",x"82",x"00", -- 0x7588
    x"39",x"34",x"10",x"0D",x"D8",x"10",x"27",x"BE", -- 0x7590
    x"B1",x"9E",x"D9",x"A6",x"80",x"9F",x"D9",x"0A", -- 0x7598
    x"D8",x"81",x"20",x"27",x"EE",x"35",x"90",x"81", -- 0x75A0
    x"3D",x"26",x"0B",x"34",x"60",x"8D",x"62",x"BD", -- 0x75A8
    x"B3",x"E9",x"DD",x"D3",x"35",x"E0",x"BD",x"F6", -- 0x75B0
    x"08",x"10",x"25",x"BE",x"8D",x"0F",x"D3",x"0F", -- 0x75B8
    x"D4",x"80",x"30",x"97",x"D7",x"DC",x"D3",x"8D", -- 0x75C0
    x"34",x"DB",x"D7",x"89",x"00",x"DD",x"D3",x"96", -- 0x75C8
    x"E6",x"81",x"02",x"2E",x"05",x"CC",x"01",x"3F", -- 0x75D0
    x"20",x"03",x"CC",x"02",x"7F",x"10",x"93",x"D3", -- 0x75D8
    x"10",x"2D",x"BE",x"66",x"DC",x"D3",x"0D",x"D8", -- 0x75E0
    x"27",x"10",x"BD",x"F5",x"91",x"BD",x"F6",x"08", -- 0x75E8
    x"24",x"CF",x"0C",x"D8",x"9E",x"D9",x"30",x"1F", -- 0x75F0
    x"9F",x"D9",x"DC",x"D3",x"39",x"58",x"49",x"34", -- 0x75F8
    x"06",x"58",x"49",x"58",x"49",x"E3",x"E1",x"39", -- 0x7600
    x"81",x"30",x"25",x"04",x"80",x"3A",x"80",x"C6", -- 0x7608
    x"39",x"9E",x"D9",x"34",x"10",x"BD",x"F5",x"91", -- 0x7610
    x"BD",x"B3",x"A2",x"10",x"25",x"BE",x"2B",x"BD", -- 0x7618
    x"F5",x"91",x"81",x"3B",x"26",x"F9",x"35",x"10", -- 0x7620
    x"DE",x"A6",x"34",x"40",x"9F",x"A6",x"BD",x"B2", -- 0x7628
    x"84",x"35",x"10",x"9F",x"A6",x"39",x"0F",x"E6", -- 0x7630
    x"10",x"21",x"09",x"C4",x"81",x"00",x"27",x"0F", -- 0x7638
    x"BD",x"B7",x"0B",x"C1",x"20",x"27",x"0B",x"C1", -- 0x7640
    x"28",x"27",x"11",x"C1",x"50",x"27",x"2A",x"7E", -- 0x7648
    x"B4",x"4A",x"4F",x"97",x"E7",x"BD",x"A9",x"28", -- 0x7650
    x"17",x"E9",x"BE",x"39",x"86",x"01",x"97",x"E7", -- 0x7658
    x"17",x"01",x"0F",x"86",x"28",x"C6",x"18",x"FD", -- 0x7660
    x"FE",x"04",x"CC",x"27",x"80",x"FD",x"FE",x"06", -- 0x7668
    x"8D",x"1A",x"17",x"01",x"03",x"17",x"E9",x"A1", -- 0x7670
    x"39",x"86",x"02",x"97",x"E7",x"17",x"00",x"F2", -- 0x7678
    x"86",x"50",x"C6",x"18",x"FD",x"FE",x"04",x"CC", -- 0x7680
    x"2F",x"00",x"20",x"E1",x"8E",x"20",x"00",x"10", -- 0x7688
    x"21",x"09",x"6D",x"BF",x"FE",x"00",x"86",x"20", -- 0x7690
    x"F6",x"FE",x"08",x"ED",x"81",x"BC",x"FE",x"06", -- 0x7698
    x"25",x"F9",x"8E",x"20",x"00",x"4F",x"B7",x"FE", -- 0x76A0
    x"02",x"B7",x"FE",x"03",x"39",x"35",x"01",x"10", -- 0x76A8
    x"21",x"09",x"4D",x"27",x"2B",x"BD",x"B7",x"0B", -- 0x76B0
    x"5D",x"27",x"25",x"C1",x"08",x"22",x"28",x"5A", -- 0x76B8
    x"31",x"8D",x"EF",x"B4",x"A6",x"A5",x"B7",x"FF", -- 0x76C0
    x"9A",x"17",x"00",x"9A",x"F7",x"FE",x"08",x"86", -- 0x76C8
    x"20",x"17",x"00",x"9E",x"8E",x"20",x"00",x"BF", -- 0x76D0
    x"FE",x"00",x"8D",x"BF",x"17",x"00",x"99",x"39", -- 0x76D8
    x"17",x"00",x"8F",x"8D",x"A7",x"20",x"F5",x"7F", -- 0x76E0
    x"FE",x"08",x"B6",x"E6",x"78",x"B7",x"FF",x"9A", -- 0x76E8
    x"8D",x"74",x"C1",x"64",x"27",x"3A",x"8D",x"7A", -- 0x76F0
    x"8D",x"92",x"8D",x"7C",x"8E",x"F7",x"01",x"7E", -- 0x76F8
    x"B9",x"9C",x"4D",x"69",x"63",x"72",x"6F",x"77", -- 0x7700
    x"61",x"72",x"65",x"20",x"53",x"79",x"73",x"74", -- 0x7708
    x"65",x"6D",x"73",x"20",x"43",x"6F",x"72",x"70", -- 0x7710
    x"2E",x"0D",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7718
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7720
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7728
    x"8D",x"40",x"17",x"FF",x"57",x"8D",x"41",x"8E", -- 0x7730
    x"F7",x"1A",x"BD",x"B9",x"9C",x"34",x"10",x"30", -- 0x7738
    x"8D",x"FF",x"B1",x"86",x"12",x"A7",x"80",x"A7", -- 0x7740
    x"84",x"30",x"8D",x"FF",x"CE",x"A7",x"80",x"8C", -- 0x7748
    x"F7",x"4D",x"25",x"F9",x"35",x"10",x"39",x"0D", -- 0x7750
    x"E7",x"26",x"06",x"BD",x"A9",x"28",x"7E",x"A3", -- 0x7758
    x"90",x"17",x"FF",x"7C",x"20",x"F8",x"34",x"20", -- 0x7760
    x"31",x"8D",x"E8",x"CF",x"A7",x"23",x"A7",x"2C", -- 0x7768
    x"35",x"A0",x"1A",x"50",x"17",x"E9",x"3E",x"39", -- 0x7770
    x"17",x"E9",x"1C",x"1C",x"AF",x"39",x"8D",x"07", -- 0x7778
    x"BD",x"A1",x"CB",x"27",x"F9",x"35",x"94",x"0A", -- 0x7780
    x"94",x"26",x"1D",x"C6",x"0B",x"D7",x"94",x"8D", -- 0x7788
    x"E1",x"BE",x"FE",x"00",x"A6",x"01",x"85",x"40", -- 0x7790
    x"27",x"05",x"B6",x"FE",x"08",x"20",x"05",x"B6", -- 0x7798
    x"FE",x"08",x"8A",x"40",x"A7",x"01",x"8D",x"D0", -- 0x77A0
    x"8E",x"04",x"5E",x"7E",x"A7",x"D3",x"8D",x"C2", -- 0x77A8
    x"10",x"21",x"08",x"4C",x"BE",x"FE",x"00",x"81", -- 0x77B0
    x"08",x"26",x"09",x"8C",x"20",x"00",x"27",x"1E", -- 0x77B8
    x"8D",x"20",x"20",x"1A",x"81",x"0D",x"26",x"04", -- 0x77C0
    x"8D",x"5D",x"20",x"0B",x"81",x"20",x"25",x"0E", -- 0x77C8
    x"F6",x"FE",x"08",x"ED",x"84",x"8D",x"30",x"BC", -- 0x77D0
    x"FE",x"06",x"25",x"02",x"8D",x"76",x"8D",x"98", -- 0x77D8
    x"35",x"96",x"34",x"06",x"86",x"20",x"F6",x"FE", -- 0x77E0
    x"08",x"ED",x"84",x"CA",x"40",x"ED",x"1E",x"30", -- 0x77E8
    x"1E",x"BF",x"FE",x"00",x"FC",x"FE",x"02",x"4A", -- 0x77F0
    x"2A",x"08",x"5A",x"F7",x"FE",x"03",x"B6",x"FE", -- 0x77F8
    x"04",x"4A",x"B7",x"FE",x"02",x"35",x"86",x"34", -- 0x7800
    x"06",x"86",x"20",x"F6",x"FE",x"08",x"CA",x"40", -- 0x7808
    x"30",x"02",x"ED",x"84",x"BF",x"FE",x"00",x"FC", -- 0x7810
    x"FE",x"02",x"4C",x"B1",x"FE",x"04",x"25",x"E2", -- 0x7818
    x"5C",x"F7",x"FE",x"03",x"4F",x"20",x"DB",x"34", -- 0x7820
    x"06",x"86",x"20",x"F6",x"FE",x"08",x"ED",x"81", -- 0x7828
    x"34",x"02",x"B6",x"FE",x"02",x"4C",x"B7",x"FE", -- 0x7830
    x"02",x"B1",x"FE",x"04",x"35",x"02",x"25",x"EE", -- 0x7838
    x"BF",x"FE",x"00",x"7F",x"FE",x"02",x"7C",x"FE", -- 0x7840
    x"03",x"86",x"20",x"F6",x"FE",x"08",x"CA",x"40", -- 0x7848
    x"ED",x"84",x"35",x"86",x"34",x"06",x"8E",x"20", -- 0x7850
    x"00",x"B6",x"FE",x"04",x"81",x"28",x"26",x"0E", -- 0x7858
    x"EC",x"88",x"50",x"ED",x"81",x"8C",x"27",x"30", -- 0x7860
    x"25",x"F6",x"8D",x"0F",x"35",x"86",x"EC",x"89", -- 0x7868
    x"00",x"A0",x"ED",x"81",x"8C",x"2E",x"60",x"25", -- 0x7870
    x"F5",x"20",x"EF",x"7F",x"FE",x"02",x"86",x"17", -- 0x7878
    x"B7",x"FE",x"03",x"86",x"20",x"F6",x"FE",x"08", -- 0x7880
    x"34",x"10",x"ED",x"81",x"BC",x"FE",x"06",x"26", -- 0x7888
    x"F9",x"7F",x"FE",x"02",x"35",x"10",x"86",x"20", -- 0x7890
    x"F6",x"FE",x"08",x"CA",x"40",x"ED",x"84",x"BF", -- 0x7898
    x"FE",x"00",x"39",x"0D",x"6F",x"26",x"04",x"0D", -- 0x78A0
    x"E7",x"26",x"06",x"BD",x"A3",x"5F",x"7E",x"B9", -- 0x78A8
    x"5F",x"17",x"FE",x"BE",x"7D",x"FE",x"02",x"34", -- 0x78B0
    x"01",x"17",x"FE",x"BC",x"35",x"01",x"10",x"26", -- 0x78B8
    x"C0",x"96",x"39",x"0D",x"E7",x"26",x"06",x"BD", -- 0x78C0
    x"A5",x"54",x"7E",x"B9",x"05",x"C6",x"4E",x"7E", -- 0x78C8
    x"AC",x"46",x"D6",x"E7",x"10",x"21",x"07",x"28", -- 0x78D0
    x"27",x"F3",x"34",x"04",x"BD",x"E7",x"B2",x"96", -- 0x78D8
    x"2C",x"35",x"04",x"C1",x"01",x"26",x"04",x"81", -- 0x78E0
    x"28",x"20",x"02",x"81",x"50",x"10",x"24",x"BB", -- 0x78E8
    x"59",x"D6",x"C0",x"C1",x"18",x"24",x"F6",x"34", -- 0x78F0
    x"06",x"17",x"FE",x"76",x"FD",x"FE",x"02",x"BE", -- 0x78F8
    x"FE",x"00",x"B6",x"FE",x"08",x"A7",x"01",x"B6", -- 0x7900
    x"FE",x"04",x"48",x"3D",x"8E",x"20",x"00",x"30", -- 0x7908
    x"8B",x"35",x"06",x"48",x"1F",x"89",x"3A",x"B6", -- 0x7910
    x"FE",x"08",x"8A",x"40",x"A7",x"01",x"BF",x"FE", -- 0x7918
    x"00",x"17",x"FE",x"54",x"39",x"0D",x"E7",x"10", -- 0x7920
    x"21",x"06",x"D5",x"27",x"A0",x"17",x"FE",x"42", -- 0x7928
    x"BE",x"FE",x"00",x"EC",x"84",x"DD",x"CB",x"FC", -- 0x7930
    x"FE",x"02",x"DD",x"CD",x"17",x"FE",x"39",x"BD", -- 0x7938
    x"B3",x"57",x"9F",x"3B",x"BD",x"B2",x"6D",x"C6", -- 0x7940
    x"01",x"BD",x"B5",x"6D",x"96",x"CB",x"BD",x"B5", -- 0x7948
    x"11",x"A7",x"84",x"BD",x"B5",x"4C",x"9E",x"3B", -- 0x7950
    x"6D",x"1F",x"10",x"2A",x"B7",x"F3",x"10",x"9E", -- 0x7958
    x"52",x"C6",x"05",x"A6",x"A0",x"A7",x"80",x"5A", -- 0x7960
    x"26",x"F9",x"9E",x"0B",x"30",x"1B",x"9F",x"0B", -- 0x7968
    x"BD",x"B3",x"57",x"9F",x"3B",x"BD",x"B2",x"6D", -- 0x7970
    x"4F",x"D6",x"CC",x"BD",x"B4",x"F4",x"9E",x"3B", -- 0x7978
    x"6D",x"1F",x"10",x"2B",x"B7",x"CB",x"BD",x"BC", -- 0x7980
    x"35",x"BD",x"B3",x"57",x"9F",x"3B",x"BD",x"B2", -- 0x7988
    x"6D",x"4F",x"D6",x"CD",x"BD",x"B4",x"F4",x"9E", -- 0x7990
    x"3B",x"6D",x"1F",x"10",x"2B",x"B7",x"B2",x"BD", -- 0x7998
    x"BC",x"35",x"BD",x"B3",x"57",x"9F",x"3B",x"4F", -- 0x79A0
    x"D6",x"CE",x"BD",x"B4",x"F4",x"9E",x"3B",x"6D", -- 0x79A8
    x"1F",x"10",x"2B",x"B7",x"9C",x"BD",x"BC",x"35", -- 0x79B0
    x"39",x"BD",x"B7",x"0B",x"10",x"21",x"06",x"40", -- 0x79B8
    x"C1",x"08",x"10",x"24",x"BA",x"84",x"58",x"58", -- 0x79C0
    x"58",x"34",x"04",x"9D",x"A5",x"BD",x"B2",x"6D", -- 0x79C8
    x"BD",x"B7",x"0B",x"C1",x"08",x"10",x"24",x"BA", -- 0x79D0
    x"71",x"EA",x"E4",x"32",x"61",x"C4",x"3F",x"34", -- 0x79D8
    x"04",x"9D",x"A5",x"27",x"21",x"BD",x"B2",x"6D", -- 0x79E0
    x"81",x"42",x"26",x"0A",x"35",x"04",x"CA",x"80", -- 0x79E8
    x"34",x"04",x"9D",x"9F",x"20",x"ED",x"81",x"55", -- 0x79F0
    x"10",x"26",x"BA",x"4E",x"35",x"04",x"CA",x"40", -- 0x79F8
    x"34",x"04",x"9D",x"9F",x"20",x"DD",x"35",x"04", -- 0x7A00
    x"F7",x"FE",x"08",x"39",x"00",x"00",x"00",x"00", -- 0x7A08
    x"38",x"44",x"40",x"40",x"40",x"44",x"38",x"10", -- 0x7A10
    x"44",x"00",x"44",x"44",x"44",x"4C",x"34",x"00", -- 0x7A18
    x"08",x"10",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7A20
    x"10",x"28",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7A28
    x"28",x"00",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7A30
    x"20",x"10",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7A38
    x"10",x"00",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7A40
    x"00",x"00",x"38",x"44",x"40",x"44",x"38",x"10", -- 0x7A48
    x"10",x"28",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7A50
    x"28",x"00",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7A58
    x"20",x"10",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7A60
    x"28",x"00",x"30",x"10",x"10",x"10",x"38",x"00", -- 0x7A68
    x"10",x"28",x"00",x"30",x"10",x"10",x"38",x"00", -- 0x7A70
    x"00",x"18",x"24",x"38",x"24",x"24",x"38",x"40", -- 0x7A78
    x"44",x"10",x"28",x"44",x"7C",x"44",x"44",x"00", -- 0x7A80
    x"10",x"10",x"28",x"44",x"7C",x"44",x"44",x"00", -- 0x7A88
    x"08",x"10",x"38",x"44",x"44",x"44",x"38",x"00", -- 0x7A90
    x"00",x"00",x"68",x"14",x"3C",x"50",x"3C",x"00", -- 0x7A98
    x"3C",x"50",x"50",x"78",x"50",x"50",x"5C",x"00", -- 0x7AA0
    x"10",x"28",x"38",x"44",x"44",x"44",x"38",x"00", -- 0x7AA8
    x"28",x"00",x"38",x"44",x"44",x"44",x"38",x"00", -- 0x7AB0
    x"00",x"00",x"38",x"4C",x"54",x"64",x"38",x"00", -- 0x7AB8
    x"10",x"28",x"00",x"44",x"44",x"4C",x"34",x"00", -- 0x7AC0
    x"20",x"10",x"44",x"44",x"44",x"4C",x"34",x"00", -- 0x7AC8
    x"38",x"4C",x"54",x"54",x"54",x"64",x"38",x"00", -- 0x7AD0
    x"44",x"38",x"44",x"44",x"44",x"44",x"38",x"00", -- 0x7AD8
    x"28",x"44",x"44",x"44",x"44",x"44",x"38",x"00", -- 0x7AE0
    x"38",x"40",x"38",x"44",x"38",x"04",x"38",x"00", -- 0x7AE8
    x"08",x"14",x"10",x"38",x"10",x"50",x"3C",x"00", -- 0x7AF0
    x"10",x"10",x"7C",x"10",x"10",x"00",x"7C",x"00", -- 0x7AF8
    x"10",x"28",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x7B00
    x"08",x"14",x"10",x"38",x"10",x"10",x"20",x"40", -- 0x7B08
    x"00",x"10",x"18",x"1C",x"1C",x"18",x"10",x"00", -- 0x7B10
    x"00",x"08",x"18",x"38",x"38",x"18",x"08",x"00", -- 0x7B18
    x"00",x"00",x"00",x"7E",x"3C",x"18",x"00",x"00", -- 0x7B20
    x"00",x"00",x"18",x"3C",x"7E",x"00",x"00",x"00", -- 0x7B28
    x"00",x"FF",x"00",x"FF",x"FF",x"00",x"FF",x"00", -- 0x7B30
    x"00",x"00",x"30",x"3C",x"14",x"1C",x"00",x"00", -- 0x7B38
    x"00",x"7E",x"42",x"5A",x"5A",x"42",x"7E",x"00", -- 0x7B40
    x"00",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"00", -- 0x7B48
    x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00", -- 0x7B50
    x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"00",x"00", -- 0x7B58
    x"00",x"7E",x"24",x"18",x"18",x"24",x"7E",x"00", -- 0x7B60
    x"00",x"7F",x"00",x"7F",x"7F",x"00",x"7F",x"00", -- 0x7B68
    x"00",x"FE",x"00",x"FE",x"FE",x"00",x"FE",x"00", -- 0x7B70
    x"38",x"44",x"40",x"40",x"40",x"44",x"38",x"10", -- 0x7B78
    x"44",x"00",x"44",x"44",x"44",x"4C",x"34",x"00", -- 0x7B80
    x"08",x"10",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7B88
    x"10",x"28",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7B90
    x"28",x"00",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7B98
    x"20",x"10",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7BA0
    x"10",x"00",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7BA8
    x"00",x"00",x"38",x"44",x"40",x"44",x"38",x"10", -- 0x7BB0
    x"10",x"28",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7BB8
    x"28",x"00",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7BC0
    x"20",x"10",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7BC8
    x"28",x"00",x"30",x"10",x"10",x"10",x"38",x"00", -- 0x7BD0
    x"10",x"28",x"00",x"30",x"10",x"10",x"38",x"00", -- 0x7BD8
    x"00",x"18",x"24",x"38",x"24",x"24",x"38",x"40", -- 0x7BE0
    x"44",x"10",x"28",x"44",x"7C",x"44",x"44",x"00", -- 0x7BE8
    x"10",x"10",x"28",x"44",x"7C",x"44",x"44",x"00", -- 0x7BF0
    x"08",x"10",x"38",x"44",x"44",x"44",x"38",x"00", -- 0x7BF8
    x"00",x"00",x"68",x"14",x"3C",x"50",x"3C",x"00", -- 0x7C00
    x"3C",x"50",x"50",x"78",x"50",x"50",x"5C",x"00", -- 0x7C08
    x"10",x"28",x"38",x"44",x"44",x"44",x"38",x"00", -- 0x7C10
    x"28",x"00",x"38",x"44",x"44",x"44",x"38",x"00", -- 0x7C18
    x"00",x"00",x"38",x"4C",x"54",x"64",x"38",x"00", -- 0x7C20
    x"10",x"28",x"00",x"44",x"44",x"4C",x"34",x"00", -- 0x7C28
    x"20",x"10",x"44",x"44",x"44",x"4C",x"34",x"00", -- 0x7C30
    x"38",x"4C",x"54",x"54",x"54",x"64",x"38",x"00", -- 0x7C38
    x"44",x"38",x"44",x"44",x"44",x"44",x"38",x"00", -- 0x7C40
    x"28",x"44",x"44",x"44",x"44",x"44",x"38",x"00", -- 0x7C48
    x"38",x"40",x"38",x"44",x"38",x"04",x"38",x"00", -- 0x7C50
    x"08",x"14",x"10",x"38",x"10",x"50",x"3C",x"00", -- 0x7C58
    x"10",x"10",x"7C",x"10",x"10",x"00",x"7C",x"00", -- 0x7C60
    x"10",x"28",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x7C68
    x"08",x"14",x"10",x"38",x"10",x"10",x"20",x"40", -- 0x7C70
    x"00",x"10",x"18",x"1C",x"1C",x"18",x"10",x"00", -- 0x7C78
    x"00",x"08",x"18",x"38",x"38",x"18",x"08",x"00", -- 0x7C80
    x"00",x"00",x"00",x"7E",x"3C",x"18",x"00",x"00", -- 0x7C88
    x"00",x"00",x"18",x"3C",x"7E",x"00",x"00",x"00", -- 0x7C90
    x"00",x"FF",x"00",x"FF",x"FF",x"00",x"FF",x"00", -- 0x7C98
    x"00",x"00",x"30",x"3C",x"14",x"1C",x"00",x"00", -- 0x7CA0
    x"00",x"7E",x"42",x"5A",x"5A",x"42",x"7E",x"00", -- 0x7CA8
    x"00",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"00", -- 0x7CB0
    x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00", -- 0x7CB8
    x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"00",x"00", -- 0x7CC0
    x"00",x"7E",x"24",x"18",x"18",x"24",x"7E",x"00", -- 0x7CC8
    x"00",x"7F",x"00",x"7F",x"7F",x"00",x"7F",x"00", -- 0x7CD0
    x"00",x"FE",x"00",x"FE",x"FE",x"00",x"FE",x"00", -- 0x7CD8
    x"38",x"44",x"40",x"40",x"40",x"44",x"38",x"10", -- 0x7CE0
    x"44",x"00",x"44",x"44",x"44",x"4C",x"34",x"00", -- 0x7CE8
    x"08",x"10",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7CF0
    x"10",x"28",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7CF8
    x"28",x"00",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7D00
    x"20",x"10",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7D08
    x"10",x"00",x"38",x"04",x"3C",x"44",x"3C",x"00", -- 0x7D10
    x"00",x"00",x"38",x"44",x"40",x"44",x"38",x"10", -- 0x7D18
    x"10",x"28",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7D20
    x"28",x"00",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7D28
    x"20",x"10",x"38",x"44",x"7C",x"40",x"38",x"00", -- 0x7D30
    x"28",x"00",x"30",x"10",x"10",x"10",x"38",x"00", -- 0x7D38
    x"10",x"28",x"00",x"30",x"10",x"10",x"38",x"00", -- 0x7D40
    x"00",x"18",x"24",x"38",x"24",x"24",x"38",x"40", -- 0x7D48
    x"44",x"10",x"28",x"44",x"7C",x"44",x"44",x"00", -- 0x7D50
    x"10",x"10",x"28",x"44",x"7C",x"44",x"44",x"00", -- 0x7D58
    x"08",x"10",x"38",x"44",x"44",x"44",x"38",x"00", -- 0x7D60
    x"00",x"00",x"68",x"14",x"3C",x"50",x"3C",x"00", -- 0x7D68
    x"3C",x"50",x"50",x"78",x"50",x"50",x"5C",x"00", -- 0x7D70
    x"10",x"28",x"38",x"44",x"44",x"44",x"38",x"00", -- 0x7D78
    x"28",x"00",x"38",x"44",x"44",x"44",x"38",x"00", -- 0x7D80
    x"00",x"00",x"38",x"4C",x"54",x"64",x"38",x"00", -- 0x7D88
    x"10",x"28",x"00",x"44",x"44",x"4C",x"34",x"00", -- 0x7D90
    x"20",x"10",x"44",x"44",x"44",x"4C",x"34",x"00", -- 0x7D98
    x"38",x"4C",x"54",x"54",x"54",x"64",x"38",x"00", -- 0x7DA0
    x"44",x"38",x"44",x"44",x"44",x"44",x"38",x"00", -- 0x7DA8
    x"28",x"44",x"44",x"44",x"44",x"44",x"38",x"00", -- 0x7DB0
    x"38",x"40",x"38",x"44",x"38",x"04",x"38",x"00", -- 0x7DB8
    x"08",x"14",x"10",x"38",x"10",x"50",x"3C",x"00", -- 0x7DC0
    x"10",x"10",x"7C",x"10",x"10",x"00",x"7C",x"00", -- 0x7DC8
    x"10",x"28",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x7DD0
    x"08",x"14",x"10",x"38",x"10",x"10",x"20",x"40", -- 0x7DD8
    x"00",x"10",x"18",x"1C",x"1C",x"18",x"10",x"00", -- 0x7DE0
    x"00",x"08",x"18",x"38",x"38",x"18",x"08",x"00", -- 0x7DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7DF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7DF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7E08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7E18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7E28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7E38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7E48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7E58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7E68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7E78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7E88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7E98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7EA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7EB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7EC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7ED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7EE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7F00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7F10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7F20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7F40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7F50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7F60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7F70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7F80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7F90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7FA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7FB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7FC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7FD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7FE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x7FE8
    x"00",x"00",x"FE",x"EE",x"FE",x"F1",x"FE",x"F4", -- 0x7FF0
    x"FE",x"F7",x"FE",x"FA",x"FE",x"FD",x"8C",x"1B", -- 0x7FF8
    x"44",x"4B",x"20",x"08",x"D7",x"5F",x"00",x"EA", -- 0x8000
    x"DF",x"4C",x"DF",x"00",x"8E",x"06",x"00",x"6F", -- 0x8008
    x"80",x"8C",x"09",x"89",x"26",x"F9",x"8E",x"C1", -- 0x8010
    x"09",x"CE",x"01",x"34",x"C6",x"0A",x"BD",x"A5", -- 0x8018
    x"9A",x"CC",x"B2",x"77",x"ED",x"43",x"ED",x"48", -- 0x8020
    x"6F",x"C4",x"6F",x"45",x"CC",x"CF",x"0A",x"FD", -- 0x8028
    x"01",x"2D",x"CC",x"CF",x"32",x"FD",x"01",x"32", -- 0x8030
    x"CE",x"01",x"5E",x"86",x"7E",x"B7",x"01",x"A0", -- 0x8038
    x"A7",x"C0",x"EC",x"81",x"ED",x"C1",x"8C",x"C1", -- 0x8040
    x"39",x"26",x"F0",x"8E",x"C2",x"B2",x"BF",x"01", -- 0x8048
    x"A1",x"8E",x"C8",x"B0",x"BF",x"01",x"9B",x"8E", -- 0x8050
    x"09",x"5F",x"9F",x"B0",x"CE",x"B4",x"4A",x"C6", -- 0x8058
    x"0A",x"EF",x"81",x"5A",x"26",x"FB",x"8E",x"D8", -- 0x8060
    x"A1",x"BF",x"01",x"0A",x"86",x"7E",x"B7",x"01", -- 0x8068
    x"09",x"8E",x"D8",x"AF",x"BF",x"01",x"0D",x"86", -- 0x8070
    x"13",x"B7",x"09",x"7A",x"7F",x"08",x"00",x"7F", -- 0x8078
    x"08",x"4A",x"7F",x"08",x"94",x"7F",x"08",x"DE", -- 0x8080
    x"8E",x"09",x"89",x"BF",x"09",x"48",x"30",x"89", -- 0x8088
    x"01",x"00",x"BF",x"09",x"4A",x"30",x"01",x"BF", -- 0x8090
    x"09",x"28",x"6F",x"00",x"30",x"89",x"01",x"19", -- 0x8098
    x"BF",x"09",x"2A",x"6F",x"00",x"30",x"89",x"01", -- 0x80A0
    x"19",x"BF",x"09",x"2C",x"6F",x"00",x"86",x"02", -- 0x80A8
    x"B7",x"09",x"5B",x"30",x"89",x"01",x"19",x"1F", -- 0x80B0
    x"10",x"5D",x"27",x"01",x"4C",x"85",x"01",x"27", -- 0x80B8
    x"01",x"4C",x"1F",x"89",x"CB",x"18",x"D7",x"19", -- 0x80C0
    x"BD",x"96",x"EC",x"96",x"BA",x"8B",x"06",x"97", -- 0x80C8
    x"B7",x"AD",x"9F",x"C0",x"08",x"8D",x"19",x"1C", -- 0x80D0
    x"AF",x"8E",x"C1",x"38",x"BD",x"B9",x"9C",x"8E", -- 0x80D8
    x"C0",x"E7",x"9F",x"72",x"7E",x"A0",x"E2",x"12", -- 0x80E0
    x"8D",x"06",x"BD",x"D2",x"D2",x"7E",x"80",x"C0", -- 0x80E8
    x"7F",x"09",x"82",x"7F",x"09",x"85",x"7F",x"09", -- 0x80F0
    x"86",x"7F",x"FF",x"40",x"86",x"D0",x"B7",x"FF", -- 0x80F8
    x"48",x"1E",x"88",x"1E",x"88",x"B6",x"FF",x"48", -- 0x8100
    x"39",x"14",x"C1",x"92",x"C2",x"38",x"06",x"C2", -- 0x8108
    x"19",x"C2",x"4E",x"C4",x"4B",x"C8",x"88",x"C8", -- 0x8110
    x"93",x"CC",x"1C",x"C5",x"BC",x"C8",x"48",x"C8", -- 0x8118
    x"4B",x"CA",x"E9",x"CA",x"F9",x"8E",x"90",x"CD", -- 0x8120
    x"35",x"C8",x"A9",x"C6",x"E4",x"CA",x"E4",x"C9", -- 0x8128
    x"0C",x"CE",x"D2",x"C6",x"E4",x"C2",x"65",x"CA", -- 0x8130
    x"3E",x"44",x"49",x"53",x"4B",x"20",x"45",x"58", -- 0x8138
    x"54",x"45",x"4E",x"44",x"45",x"44",x"20",x"43", -- 0x8140
    x"4F",x"4C",x"4F",x"52",x"20",x"42",x"41",x"53", -- 0x8148
    x"49",x"43",x"20",x"31",x"2E",x"31",x"0D",x"43", -- 0x8150
    x"4F",x"50",x"59",x"52",x"49",x"47",x"48",x"54", -- 0x8158
    x"20",x"28",x"43",x"29",x"20",x"31",x"39",x"38", -- 0x8160
    x"32",x"20",x"42",x"59",x"20",x"54",x"41",x"4E", -- 0x8168
    x"44",x"59",x"0D",x"55",x"4E",x"44",x"45",x"52", -- 0x8170
    x"20",x"4C",x"49",x"43",x"45",x"4E",x"53",x"45", -- 0x8178
    x"20",x"46",x"52",x"4F",x"4D",x"20",x"4D",x"49", -- 0x8180
    x"43",x"52",x"4F",x"53",x"4F",x"46",x"54",x"0D", -- 0x8188
    x"0D",x"00",x"44",x"49",x"D2",x"44",x"52",x"49", -- 0x8190
    x"56",x"C5",x"46",x"49",x"45",x"4C",x"C4",x"46", -- 0x8198
    x"49",x"4C",x"45",x"D3",x"4B",x"49",x"4C",x"CC", -- 0x81A0
    x"4C",x"4F",x"41",x"C4",x"4C",x"53",x"45",x"D4", -- 0x81A8
    x"4D",x"45",x"52",x"47",x"C5",x"52",x"45",x"4E", -- 0x81B0
    x"41",x"4D",x"C5",x"52",x"53",x"45",x"D4",x"53", -- 0x81B8
    x"41",x"56",x"C5",x"57",x"52",x"49",x"54",x"C5", -- 0x81C0
    x"56",x"45",x"52",x"49",x"46",x"D9",x"55",x"4E", -- 0x81C8
    x"4C",x"4F",x"41",x"C4",x"44",x"53",x"4B",x"49", -- 0x81D0
    x"4E",x"C9",x"42",x"41",x"43",x"4B",x"55",x"D0", -- 0x81D8
    x"43",x"4F",x"50",x"D9",x"44",x"53",x"4B",x"49", -- 0x81E0
    x"A4",x"44",x"53",x"4B",x"4F",x"A4",x"44",x"4F", -- 0x81E8
    x"D3",x"CC",x"A9",x"CE",x"C5",x"D0",x"BC",x"D1", -- 0x81F0
    x"5C",x"C6",x"EF",x"CA",x"48",x"D1",x"02",x"CA", -- 0x81F8
    x"39",x"D0",x"1B",x"D1",x"01",x"C9",x"E0",x"D0", -- 0x8200
    x"66",x"D7",x"4E",x"D2",x"33",x"D5",x"99",x"D2", -- 0x8208
    x"62",x"D3",x"B9",x"D4",x"ED",x"D5",x"62",x"D6", -- 0x8210
    x"EC",x"43",x"56",x"CE",x"46",x"52",x"45",x"C5", -- 0x8218
    x"4C",x"4F",x"C3",x"4C",x"4F",x"C6",x"4D",x"4B", -- 0x8220
    x"4E",x"A4",x"41",x"D3",x"CD",x"F4",x"CE",x"9C", -- 0x8228
    x"CE",x"10",x"CE",x"37",x"CE",x"02",x"B2",x"77", -- 0x8230
    x"81",x"E1",x"22",x"08",x"8E",x"C1",x"F1",x"80", -- 0x8238
    x"CE",x"7E",x"AD",x"D4",x"81",x"E1",x"10",x"23", -- 0x8240
    x"F0",x"2D",x"6E",x"9F",x"01",x"41",x"C1",x"4E", -- 0x8248
    x"23",x"04",x"6E",x"9F",x"01",x"46",x"C0",x"44", -- 0x8250
    x"34",x"04",x"BD",x"B2",x"62",x"35",x"04",x"8E", -- 0x8258
    x"C2",x"2C",x"7E",x"B2",x"CE",x"35",x"20",x"BD", -- 0x8260
    x"AD",x"33",x"BD",x"D2",x"D2",x"34",x"24",x"BD", -- 0x8268
    x"CA",x"E9",x"35",x"04",x"C1",x"36",x"10",x"25", -- 0x8270
    x"C6",x"76",x"32",x"62",x"BD",x"A7",x"E9",x"BD", -- 0x8278
    x"A9",x"74",x"0F",x"6F",x"BD",x"B9",x"5C",x"BD", -- 0x8280
    x"B9",x"AF",x"8E",x"C2",x"5A",x"7E",x"AC",x"60", -- 0x8288
    x"42",x"52",x"44",x"46",x"4F",x"42",x"57",x"50", -- 0x8290
    x"46",x"4E",x"46",x"53",x"41",x"45",x"46",x"4F", -- 0x8298
    x"53",x"45",x"56",x"46",x"45",x"52",x"42",x"41", -- 0x82A0
    x"53",x"20",x"20",x"20",x"44",x"41",x"54",x"42", -- 0x82A8
    x"49",x"4E",x"34",x"11",x"AE",x"63",x"8C",x"97", -- 0x82B0
    x"5F",x"26",x"04",x"81",x"23",x"27",x"02",x"35", -- 0x82B8
    x"91",x"32",x"65",x"BD",x"C8",x"2E",x"9F",x"F1", -- 0x82C0
    x"6F",x"88",x"15",x"6F",x"88",x"16",x"6F",x"88", -- 0x82C8
    x"17",x"6F",x"88",x"18",x"6F",x"06",x"A6",x"01", -- 0x82D0
    x"97",x"EB",x"9D",x"A5",x"27",x"0C",x"BD",x"B2", -- 0x82D8
    x"6D",x"BD",x"B7",x"3D",x"1F",x"10",x"9E",x"F1", -- 0x82E0
    x"ED",x"07",x"EC",x"07",x"27",x"1D",x"BD",x"C6", -- 0x82E8
    x"85",x"EC",x"09",x"AE",x"0B",x"34",x"16",x"30", -- 0x82F0
    x"5E",x"BD",x"9F",x"B5",x"34",x"60",x"A6",x"E0", -- 0x82F8
    x"26",x"09",x"35",x"10",x"35",x"04",x"8C",x"02", -- 0x8300
    x"64",x"25",x"05",x"C6",x"36",x"7E",x"AC",x"46", -- 0x8308
    x"DE",x"F1",x"AC",x"4D",x"10",x"27",x"00",x"B7", -- 0x8310
    x"34",x"14",x"A6",x"4F",x"27",x"06",x"6F",x"4F", -- 0x8318
    x"C6",x"03",x"8D",x"33",x"EC",x"61",x"BD",x"C7", -- 0x8320
    x"84",x"34",x"04",x"BD",x"C7",x"79",x"50",x"EB", -- 0x8328
    x"63",x"5C",x"E7",x"44",x"E6",x"42",x"BD",x"C7", -- 0x8330
    x"55",x"33",x"06",x"A6",x"E4",x"4C",x"30",x"C4", -- 0x8338
    x"3A",x"4A",x"27",x"37",x"E7",x"E4",x"E6",x"84", -- 0x8340
    x"C1",x"C0",x"25",x"F2",x"E6",x"E4",x"0D",x"D8", -- 0x8348
    x"26",x"14",x"C6",x"2E",x"7E",x"AC",x"46",x"30", -- 0x8350
    x"C8",x"19",x"D7",x"EA",x"9F",x"EE",x"30",x"C4", -- 0x8358
    x"BD",x"C7",x"63",x"7E",x"D6",x"F2",x"34",x"12", -- 0x8360
    x"BD",x"C7",x"BF",x"1F",x"89",x"35",x"42",x"E7", -- 0x8368
    x"C4",x"4A",x"26",x"F2",x"34",x"14",x"BD",x"C7", -- 0x8370
    x"1E",x"35",x"14",x"32",x"61",x"DE",x"F1",x"E7", -- 0x8378
    x"43",x"86",x"FF",x"A7",x"4D",x"A6",x"84",x"81", -- 0x8380
    x"C0",x"25",x"27",x"84",x"3F",x"A1",x"44",x"24", -- 0x8388
    x"21",x"96",x"D8",x"27",x"BD",x"A6",x"44",x"8A", -- 0x8390
    x"C0",x"A7",x"84",x"BD",x"C5",x"A9",x"AE",x"49", -- 0x8398
    x"8C",x"01",x"00",x"26",x"08",x"AC",x"C8",x"13", -- 0x83A0
    x"27",x"08",x"86",x"81",x"21",x"4F",x"5F",x"ED", -- 0x83A8
    x"C8",x"13",x"C6",x"02",x"AE",x"49",x"8C",x"01", -- 0x83B0
    x"00",x"26",x"0D",x"32",x"67",x"AE",x"4B",x"96", -- 0x83B8
    x"D8",x"27",x"02",x"C6",x"03",x"7E",x"C3",x"5A", -- 0x83C0
    x"BD",x"C3",x"57",x"35",x"14",x"AF",x"4D",x"34", -- 0x83C8
    x"04",x"BD",x"C7",x"55",x"30",x"06",x"E6",x"43", -- 0x83D0
    x"3A",x"A6",x"84",x"81",x"C0",x"25",x"2B",x"84", -- 0x83D8
    x"3F",x"A1",x"44",x"26",x"25",x"EC",x"C8",x"13", -- 0x83E0
    x"84",x"7F",x"34",x"06",x"4F",x"E6",x"62",x"E3", -- 0x83E8
    x"63",x"10",x"A3",x"E1",x"23",x"14",x"0D",x"D8", -- 0x83F0
    x"10",x"27",x"FF",x"56",x"10",x"83",x"01",x"00", -- 0x83F8
    x"23",x"03",x"CC",x"01",x"00",x"8A",x"80",x"ED", -- 0x8400
    x"C8",x"13",x"35",x"04",x"30",x"C8",x"19",x"3A", -- 0x8408
    x"EE",x"62",x"34",x"04",x"86",x"FF",x"E3",x"61", -- 0x8410
    x"24",x"07",x"ED",x"61",x"35",x"04",x"50",x"20", -- 0x8418
    x"08",x"E6",x"62",x"6F",x"61",x"6F",x"62",x"32", -- 0x8420
    x"61",x"96",x"D8",x"27",x"02",x"1E",x"13",x"BD", -- 0x8428
    x"A5",x"9A",x"EF",x"62",x"DE",x"F1",x"96",x"D8", -- 0x8430
    x"27",x"04",x"A7",x"4F",x"AF",x"62",x"AE",x"4D", -- 0x8438
    x"30",x"01",x"5F",x"EE",x"E4",x"10",x"26",x"FE", -- 0x8440
    x"BD",x"35",x"96",x"32",x"62",x"BD",x"B1",x"56", -- 0x8448
    x"BD",x"B6",x"A4",x"34",x"04",x"BD",x"A5",x"A2", -- 0x8450
    x"5D",x"10",x"2F",x"E1",x"A6",x"35",x"02",x"34", -- 0x8458
    x"06",x"0F",x"6F",x"BD",x"B2",x"6D",x"8E",x"C2", -- 0x8460
    x"AC",x"BD",x"C9",x"38",x"CC",x"01",x"FF",x"FD", -- 0x8468
    x"09",x"57",x"8E",x"01",x"00",x"9D",x"A5",x"27", -- 0x8470
    x"08",x"BD",x"B2",x"6D",x"BD",x"B3",x"E6",x"9E", -- 0x8478
    x"52",x"BF",x"09",x"7C",x"10",x"27",x"EF",x"C2", -- 0x8480
    x"BD",x"A5",x"C7",x"35",x"06",x"34",x"02",x"BD", -- 0x8488
    x"C7",x"49",x"10",x"26",x"E1",x"86",x"9F",x"F1", -- 0x8490
    x"BD",x"C7",x"9D",x"BD",x"C6",x"8C",x"35",x"04", -- 0x8498
    x"86",x"10",x"34",x"02",x"C1",x"49",x"26",x"1F", -- 0x84A0
    x"BD",x"C6",x"E5",x"BD",x"C8",x"07",x"BE",x"09", -- 0x84A8
    x"74",x"EC",x"0B",x"FD",x"09",x"57",x"8D",x"75", -- 0x84B0
    x"BD",x"C6",x"27",x"BD",x"C7",x"55",x"6C",x"00", -- 0x84B8
    x"9E",x"F1",x"35",x"02",x"A7",x"00",x"39",x"68", -- 0x84C0
    x"E4",x"C1",x"4F",x"26",x"1B",x"7D",x"09",x"73", -- 0x84C8
    x"27",x"0F",x"BD",x"C6",x"FC",x"B6",x"09",x"73", -- 0x84D0
    x"B7",x"09",x"77",x"BE",x"09",x"74",x"BF",x"09", -- 0x84D8
    x"78",x"BD",x"C5",x"67",x"8D",x"52",x"20",x"D3", -- 0x84E0
    x"C1",x"52",x"27",x"06",x"C1",x"44",x"10",x"26", -- 0x84E8
    x"E1",x"24",x"68",x"E4",x"FC",x"09",x"48",x"34", -- 0x84F0
    x"06",x"F3",x"09",x"7C",x"25",x"06",x"10",x"B3", -- 0x84F8
    x"09",x"4A",x"23",x"05",x"C6",x"3A",x"7E",x"AC", -- 0x8500
    x"46",x"34",x"06",x"7D",x"09",x"73",x"26",x"04", -- 0x8508
    x"8D",x"55",x"20",x"05",x"86",x"FF",x"BD",x"C8", -- 0x8510
    x"07",x"8D",x"12",x"63",x"0D",x"6C",x"08",x"35", -- 0x8518
    x"46",x"FD",x"09",x"48",x"EF",x"0B",x"FE",x"09", -- 0x8520
    x"7C",x"EF",x"09",x"20",x"8E",x"8D",x"09",x"FE", -- 0x8528
    x"09",x"74",x"EE",x"4E",x"EF",x"88",x"13",x"39", -- 0x8530
    x"9E",x"F1",x"C6",x"19",x"6F",x"80",x"5A",x"26", -- 0x8538
    x"FB",x"9E",x"F1",x"96",x"EB",x"A7",x"01",x"B6", -- 0x8540
    x"09",x"76",x"A7",x"02",x"A7",x"03",x"F6",x"09", -- 0x8548
    x"73",x"C0",x"03",x"58",x"58",x"58",x"34",x"04", -- 0x8550
    x"FC",x"09",x"74",x"83",x"06",x"00",x"86",x"08", -- 0x8558
    x"3D",x"AB",x"E0",x"A7",x"88",x"12",x"39",x"C6", -- 0x8560
    x"38",x"B6",x"09",x"77",x"10",x"27",x"E6",x"D6", -- 0x8568
    x"B7",x"09",x"73",x"97",x"ED",x"C6",x"02",x"D7", -- 0x8570
    x"EA",x"BD",x"D6",x"F2",x"BE",x"09",x"78",x"BF", -- 0x8578
    x"09",x"74",x"33",x"84",x"C6",x"20",x"6F",x"80", -- 0x8580
    x"5A",x"26",x"FB",x"8E",x"09",x"4C",x"C6",x"0B", -- 0x8588
    x"BD",x"A5",x"9A",x"FC",x"09",x"57",x"ED",x"40", -- 0x8590
    x"C6",x"21",x"BD",x"C7",x"BF",x"B7",x"09",x"76", -- 0x8598
    x"A7",x"42",x"C6",x"03",x"D7",x"EA",x"BD",x"D6", -- 0x85A0
    x"F2",x"34",x"56",x"BD",x"C7",x"55",x"6C",x"01", -- 0x85A8
    x"A6",x"01",x"B1",x"09",x"7A",x"25",x"03",x"BD", -- 0x85B0
    x"C7",x"1E",x"35",x"D6",x"96",x"6F",x"10",x"2F", -- 0x85B8
    x"C7",x"2F",x"32",x"62",x"34",x"14",x"0F",x"70", -- 0x85C0
    x"8E",x"09",x"26",x"D6",x"6F",x"58",x"AE",x"85", -- 0x85C8
    x"E6",x"84",x"C1",x"40",x"26",x"16",x"EC",x"88", -- 0x85D0
    x"15",x"10",x"A3",x"09",x"24",x"20",x"C3",x"00", -- 0x85D8
    x"01",x"ED",x"88",x"15",x"AE",x"0B",x"30",x"8B", -- 0x85E0
    x"A6",x"1F",x"35",x"94",x"E6",x"88",x"10",x"27", -- 0x85E8
    x"08",x"A6",x"88",x"11",x"6F",x"88",x"10",x"35", -- 0x85F0
    x"94",x"E6",x"88",x"17",x"27",x"04",x"03",x"70", -- 0x85F8
    x"35",x"94",x"E6",x"05",x"6C",x"05",x"6A",x"88", -- 0x8600
    x"18",x"27",x"06",x"3A",x"A6",x"88",x"19",x"35", -- 0x8608
    x"94",x"34",x"60",x"4F",x"33",x"8B",x"A6",x"C8", -- 0x8610
    x"19",x"34",x"02",x"6F",x"05",x"A6",x"01",x"97", -- 0x8618
    x"EB",x"8D",x"04",x"35",x"62",x"35",x"94",x"A6", -- 0x8620
    x"04",x"4C",x"34",x"02",x"81",x"09",x"23",x"01", -- 0x8628
    x"4F",x"A7",x"04",x"E6",x"03",x"33",x"84",x"BD", -- 0x8630
    x"C7",x"55",x"3A",x"E6",x"06",x"30",x"C4",x"C1", -- 0x8638
    x"C0",x"24",x"0A",x"35",x"02",x"80",x"0A",x"26", -- 0x8640
    x"15",x"E7",x"03",x"20",x"DC",x"C4",x"3F",x"C1", -- 0x8648
    x"09",x"23",x"05",x"C6",x"40",x"7E",x"AC",x"46", -- 0x8650
    x"E0",x"E0",x"25",x"21",x"1F",x"98",x"34",x"02", -- 0x8658
    x"8D",x"23",x"86",x"02",x"97",x"EA",x"BD",x"C7", -- 0x8660
    x"63",x"33",x"88",x"19",x"DF",x"EE",x"BD",x"D6", -- 0x8668
    x"F2",x"6F",x"88",x"18",x"E6",x"E0",x"26",x"0C", -- 0x8670
    x"EC",x"88",x"13",x"26",x"04",x"5F",x"63",x"88", -- 0x8678
    x"17",x"E7",x"88",x"18",x"39",x"EE",x"07",x"33", -- 0x8680
    x"41",x"EF",x"07",x"39",x"7F",x"09",x"73",x"7F", -- 0x8688
    x"09",x"77",x"CC",x"11",x"02",x"97",x"EC",x"D7", -- 0x8690
    x"EA",x"C6",x"03",x"D7",x"ED",x"CE",x"06",x"00", -- 0x8698
    x"DF",x"EE",x"BD",x"D6",x"F2",x"FF",x"09",x"74", -- 0x86A0
    x"31",x"C4",x"A6",x"C4",x"26",x"28",x"8D",x"29", -- 0x86A8
    x"8E",x"09",x"4C",x"A6",x"80",x"A1",x"C0",x"26", -- 0x86B0
    x"0E",x"8C",x"09",x"57",x"26",x"F5",x"F7",x"09", -- 0x86B8
    x"73",x"A6",x"42",x"B7",x"09",x"76",x"39",x"33", -- 0x86C0
    x"A8",x"20",x"11",x"83",x"07",x"00",x"26",x"D5", -- 0x86C8
    x"5C",x"C1",x"0B",x"23",x"C6",x"39",x"43",x"26", -- 0x86D0
    x"D7",x"B6",x"09",x"77",x"26",x"06",x"F7",x"09", -- 0x86D8
    x"77",x"FF",x"09",x"78",x"39",x"C6",x"34",x"7D", -- 0x86E0
    x"09",x"73",x"26",x"F8",x"7E",x"AC",x"46",x"BD", -- 0x86E8
    x"C9",x"35",x"BD",x"A5",x"C7",x"BD",x"C7",x"9D", -- 0x86F0
    x"8D",x"92",x"8D",x"E9",x"86",x"FF",x"BD",x"C8", -- 0x86F8
    x"07",x"BE",x"09",x"74",x"6F",x"84",x"C6",x"03", -- 0x8700
    x"D7",x"EA",x"BD",x"D6",x"F2",x"E6",x"0D",x"8D", -- 0x8708
    x"44",x"30",x"06",x"3A",x"E6",x"84",x"86",x"FF", -- 0x8710
    x"A7",x"84",x"C1",x"C0",x"25",x"F1",x"CE",x"06", -- 0x8718
    x"00",x"DF",x"EE",x"CC",x"11",x"03",x"97",x"EC", -- 0x8720
    x"D7",x"EA",x"C6",x"02",x"D7",x"ED",x"8D",x"25", -- 0x8728
    x"6F",x"01",x"30",x"06",x"C6",x"44",x"BD",x"A5", -- 0x8730
    x"9A",x"6F",x"C0",x"11",x"83",x"07",x"00",x"26", -- 0x8738
    x"F8",x"7E",x"D6",x"F2",x"34",x"04",x"D6",x"6F", -- 0x8740
    x"8C",x"34",x"04",x"58",x"8E",x"09",x"26",x"AE", -- 0x8748
    x"85",x"E6",x"00",x"35",x"84",x"34",x"06",x"96", -- 0x8750
    x"EB",x"C6",x"4A",x"3D",x"8E",x"08",x"00",x"30", -- 0x8758
    x"8B",x"35",x"86",x"E6",x"03",x"54",x"D7",x"EC", -- 0x8760
    x"C1",x"11",x"25",x"02",x"0C",x"EC",x"58",x"50", -- 0x8768
    x"EB",x"03",x"8D",x"05",x"EB",x"04",x"D7",x"ED", -- 0x8770
    x"39",x"34",x"06",x"58",x"49",x"58",x"49",x"58", -- 0x8778
    x"49",x"E3",x"E1",x"39",x"6F",x"E2",x"6C",x"E4", -- 0x8780
    x"83",x"00",x"5A",x"2A",x"F9",x"A6",x"E4",x"E7", -- 0x8788
    x"E4",x"C6",x"0A",x"3D",x"35",x"02",x"5A",x"8B", -- 0x8790
    x"09",x"2B",x"FB",x"4F",x"39",x"8D",x"B6",x"6D", -- 0x8798
    x"00",x"26",x"F9",x"6F",x"01",x"33",x"06",x"8E", -- 0x87A0
    x"06",x"00",x"9F",x"EE",x"CC",x"11",x"02",x"97", -- 0x87A8
    x"EC",x"D7",x"EA",x"C6",x"02",x"D7",x"ED",x"BD", -- 0x87B0
    x"D6",x"F2",x"C6",x"44",x"7E",x"A5",x"9A",x"8D", -- 0x87B8
    x"94",x"30",x"06",x"4F",x"C4",x"FE",x"6F",x"E2", -- 0x87C0
    x"63",x"85",x"27",x"31",x"63",x"85",x"4C",x"81", -- 0x87C8
    x"44",x"24",x"25",x"5C",x"C5",x"01",x"26",x"F0", -- 0x87D0
    x"34",x"06",x"C0",x"02",x"63",x"62",x"26",x"0C", -- 0x87D8
    x"E0",x"E0",x"2A",x"04",x"E6",x"E4",x"63",x"61", -- 0x87E0
    x"32",x"61",x"20",x"DC",x"EB",x"E0",x"C1",x"44", -- 0x87E8
    x"25",x"F6",x"E6",x"E4",x"C0",x"04",x"20",x"EE", -- 0x87F0
    x"C6",x"38",x"7E",x"AC",x"46",x"32",x"61",x"1F", -- 0x87F8
    x"98",x"3A",x"C6",x"C0",x"E7",x"84",x"39",x"34", -- 0x8800
    x"02",x"F6",x"09",x"5B",x"5C",x"BD",x"C7",x"49", -- 0x8808
    x"27",x"17",x"96",x"EB",x"A1",x"01",x"26",x"11", -- 0x8810
    x"FE",x"09",x"74",x"A6",x"4D",x"A1",x"02",x"26", -- 0x8818
    x"08",x"A6",x"00",x"A1",x"E4",x"10",x"26",x"DD", -- 0x8820
    x"F3",x"5A",x"26",x"E1",x"35",x"82",x"BD",x"A5", -- 0x8828
    x"A5",x"0F",x"6F",x"5D",x"10",x"2F",x"EC",x"12", -- 0x8830
    x"BD",x"C7",x"49",x"A6",x"00",x"10",x"27",x"DB", -- 0x8838
    x"BA",x"81",x"40",x"27",x"C1",x"7E",x"A6",x"16", -- 0x8840
    x"86",x"10",x"8C",x"86",x"20",x"0D",x"6F",x"2F", -- 0x8848
    x"B5",x"AF",x"E4",x"BD",x"C7",x"44",x"34",x"06", -- 0x8850
    x"A6",x"00",x"10",x"27",x"DB",x"9D",x"81",x"40", -- 0x8858
    x"27",x"06",x"A1",x"E4",x"26",x"DF",x"35",x"96", -- 0x8860
    x"AE",x"64",x"8C",x"B0",x"0C",x"26",x"F7",x"BD", -- 0x8868
    x"B2",x"6D",x"81",x"22",x"26",x"0B",x"BD",x"B2", -- 0x8870
    x"44",x"BD",x"B6",x"57",x"C6",x"3B",x"BD",x"B2", -- 0x8878
    x"6F",x"8E",x"B0",x"1E",x"AF",x"64",x"35",x"96", -- 0x8880
    x"2F",x"25",x"F1",x"09",x"5B",x"10",x"22",x"DD", -- 0x8888
    x"8E",x"35",x"90",x"0D",x"6F",x"2F",x"18",x"32", -- 0x8890
    x"62",x"34",x"16",x"0F",x"6E",x"BD",x"C7",x"44", -- 0x8898
    x"E6",x"06",x"4F",x"8E",x"10",x"00",x"7E",x"A3", -- 0x88A0
    x"7C",x"0D",x"6F",x"2F",x"02",x"32",x"62",x"39", -- 0x88A8
    x"32",x"62",x"1C",x"AF",x"7F",x"FF",x"02",x"B6", -- 0x88B0
    x"FF",x"00",x"43",x"84",x"7F",x"27",x"03",x"BD", -- 0x88B8
    x"AD",x"EB",x"9E",x"A6",x"9F",x"2F",x"A6",x"80", -- 0x88C0
    x"27",x"07",x"81",x"3A",x"27",x"25",x"7E",x"B2", -- 0x88C8
    x"77",x"A6",x"81",x"97",x"00",x"26",x"03",x"7E", -- 0x88D0
    x"AE",x"15",x"EC",x"80",x"DD",x"68",x"9F",x"A6", -- 0x88D8
    x"96",x"AF",x"27",x"0F",x"86",x"5B",x"BD",x"A2", -- 0x88E0
    x"82",x"96",x"68",x"BD",x"BD",x"CC",x"86",x"5D", -- 0x88E8
    x"BD",x"A2",x"82",x"9D",x"9F",x"1F",x"A9",x"81", -- 0x88F0
    x"98",x"26",x"03",x"7E",x"83",x"16",x"81",x"97", -- 0x88F8
    x"26",x"03",x"7E",x"83",x"11",x"1F",x"9A",x"BD", -- 0x8900
    x"AD",x"C6",x"20",x"A6",x"32",x"62",x"96",x"6F", -- 0x8908
    x"34",x"02",x"BD",x"A5",x"AE",x"BD",x"A3",x"ED", -- 0x8910
    x"0D",x"6F",x"10",x"2F",x"DC",x"BC",x"BD",x"C7", -- 0x8918
    x"44",x"E6",x"00",x"C1",x"40",x"10",x"27",x"DC", -- 0x8920
    x"ED",x"5F",x"A6",x"88",x"10",x"26",x"03",x"E6", -- 0x8928
    x"88",x"17",x"7E",x"A5",x"E4",x"8E",x"C2",x"A9", -- 0x8930
    x"6F",x"E2",x"B6",x"09",x"5A",x"97",x"EB",x"CE", -- 0x8938
    x"09",x"4C",x"CC",x"20",x"08",x"A7",x"C0",x"5A", -- 0x8940
    x"26",x"FB",x"C6",x"03",x"BD",x"A5",x"9A",x"BD", -- 0x8948
    x"87",x"48",x"33",x"84",x"C1",x"02",x"25",x"12", -- 0x8950
    x"A6",x"41",x"81",x"3A",x"26",x"0C",x"A6",x"C4", -- 0x8958
    x"81",x"30",x"25",x"06",x"81",x"33",x"22",x"02", -- 0x8960
    x"8D",x"33",x"8E",x"09",x"4C",x"5C",x"5A",x"26", -- 0x8968
    x"0C",x"32",x"61",x"8C",x"09",x"4C",x"26",x"67", -- 0x8970
    x"C6",x"3E",x"7E",x"AC",x"46",x"A6",x"C0",x"81", -- 0x8978
    x"2E",x"27",x"2D",x"81",x"2F",x"27",x"29",x"81", -- 0x8980
    x"3A",x"27",x"09",x"8C",x"09",x"54",x"27",x"E8", -- 0x8988
    x"8D",x"3E",x"20",x"DA",x"8D",x"DD",x"8D",x"05", -- 0x8990
    x"5D",x"26",x"DD",x"35",x"82",x"63",x"62",x"27", -- 0x8998
    x"D7",x"A6",x"C1",x"C0",x"02",x"80",x"30",x"25", -- 0x89A0
    x"CF",x"81",x"03",x"22",x"CB",x"97",x"EB",x"39", -- 0x89A8
    x"8D",x"C1",x"8E",x"09",x"57",x"86",x"20",x"A7", -- 0x89B0
    x"82",x"8C",x"09",x"54",x"26",x"F9",x"5A",x"27", -- 0x89B8
    x"DA",x"A6",x"C0",x"81",x"3A",x"27",x"CD",x"8C", -- 0x89C0
    x"09",x"57",x"27",x"AC",x"8D",x"02",x"20",x"EE", -- 0x89C8
    x"A7",x"80",x"27",x"A4",x"81",x"2E",x"27",x"A0", -- 0x89D0
    x"81",x"2F",x"27",x"9C",x"4C",x"27",x"99",x"39", -- 0x89D8
    x"81",x"4D",x"10",x"27",x"05",x"82",x"8D",x"4B", -- 0x89E0
    x"9E",x"8A",x"BF",x"09",x"57",x"9D",x"A5",x"27", -- 0x89E8
    x"21",x"BD",x"B2",x"6D",x"C6",x"41",x"BD",x"B2", -- 0x89F0
    x"6F",x"26",x"E4",x"73",x"09",x"58",x"8D",x"04", -- 0x89F8
    x"4F",x"7E",x"B7",x"64",x"86",x"4F",x"8C",x"86", -- 0x8A00
    x"49",x"F6",x"09",x"5B",x"5C",x"D7",x"6F",x"7E", -- 0x8A08
    x"C4",x"8D",x"8D",x"F0",x"86",x"FF",x"BD",x"CC", -- 0x8A10
    x"24",x"DC",x"1B",x"93",x"19",x"BD",x"CC",x"24", -- 0x8A18
    x"1F",x"98",x"BD",x"CC",x"24",x"9E",x"19",x"A6", -- 0x8A20
    x"80",x"BD",x"CC",x"24",x"9C",x"1B",x"26",x"F7", -- 0x8A28
    x"7E",x"A4",x"2D",x"8E",x"C2",x"A6",x"7E",x"C9", -- 0x8A30
    x"38",x"4F",x"C6",x"FF",x"20",x"12",x"81",x"22", -- 0x8A38
    x"10",x"26",x"B8",x"58",x"86",x"02",x"20",x"07", -- 0x8A40
    x"81",x"4D",x"10",x"27",x"05",x"73",x"4F",x"5F", -- 0x8A48
    x"B7",x"09",x"59",x"F7",x"09",x"5E",x"8D",x"DB", -- 0x8A50
    x"9D",x"A5",x"27",x"10",x"BD",x"B2",x"6D",x"C6", -- 0x8A58
    x"52",x"BD",x"B2",x"6F",x"BD",x"A5",x"C7",x"86", -- 0x8A60
    x"03",x"B7",x"09",x"59",x"8D",x"99",x"B6",x"09", -- 0x8A68
    x"58",x"27",x"0B",x"7D",x"09",x"5E",x"26",x"03", -- 0x8A70
    x"BD",x"AD",x"19",x"7E",x"AC",x"7C",x"B6",x"09", -- 0x8A78
    x"57",x"BA",x"09",x"5E",x"10",x"26",x"DB",x"8E", -- 0x8A80
    x"BD",x"AD",x"19",x"73",x"09",x"5D",x"BD",x"CD", -- 0x8A88
    x"BC",x"BD",x"CD",x"BC",x"34",x"02",x"BD",x"CD", -- 0x8A90
    x"BC",x"1F",x"89",x"35",x"02",x"D3",x"19",x"BD", -- 0x8A98
    x"AC",x"37",x"9E",x"19",x"BD",x"C5",x"C4",x"D6", -- 0x8AA0
    x"70",x"26",x"04",x"A7",x"80",x"20",x"F5",x"7F", -- 0x8AA8
    x"09",x"5D",x"9F",x"1B",x"C6",x"03",x"A6",x"82", -- 0x8AB0
    x"26",x"03",x"5A",x"26",x"F9",x"9E",x"1B",x"9F", -- 0x8AB8
    x"1B",x"6F",x"80",x"5A",x"2A",x"F9",x"BD",x"A4", -- 0x8AC0
    x"2D",x"BD",x"AD",x"21",x"BD",x"82",x"9C",x"BD", -- 0x8AC8
    x"AC",x"EF",x"77",x"09",x"59",x"25",x"03",x"BD", -- 0x8AD0
    x"A4",x"26",x"77",x"09",x"59",x"10",x"25",x"E2", -- 0x8AD8
    x"BD",x"7E",x"AC",x"73",x"0D",x"6F",x"2E",x"DE", -- 0x8AE0
    x"39",x"F6",x"09",x"5B",x"5C",x"34",x"04",x"D7", -- 0x8AE8
    x"6F",x"8D",x"0E",x"35",x"04",x"5A",x"26",x"F5", -- 0x8AF0
    x"39",x"0D",x"6F",x"10",x"2F",x"B7",x"87",x"32", -- 0x8AF8
    x"62",x"BD",x"C7",x"44",x"0F",x"6F",x"9F",x"F1", -- 0x8B00
    x"A6",x"00",x"27",x"EC",x"34",x"02",x"6F",x"00", -- 0x8B08
    x"E6",x"01",x"D7",x"EB",x"81",x"20",x"26",x"19", -- 0x8B10
    x"E6",x"88",x"18",x"86",x"80",x"AA",x"05",x"ED", -- 0x8B18
    x"88",x"13",x"6C",x"04",x"E6",x"03",x"BD",x"C7", -- 0x8B20
    x"55",x"A7",x"01",x"3A",x"6C",x"06",x"7E",x"CB", -- 0x8B28
    x"C3",x"81",x"40",x"26",x"F9",x"EC",x"09",x"AE", -- 0x8B30
    x"0B",x"31",x"8B",x"34",x"36",x"31",x"E4",x"DE", -- 0x8B38
    x"1B",x"11",x"93",x"1D",x"27",x"0E",x"A6",x"41", -- 0x8B40
    x"33",x"42",x"2A",x"02",x"8D",x"28",x"33",x"45", -- 0x8B48
    x"20",x"EF",x"35",x"40",x"11",x"93",x"1F",x"27", -- 0x8B50
    x"3A",x"1F",x"30",x"E3",x"42",x"34",x"06",x"A6", -- 0x8B58
    x"41",x"2A",x"EF",x"E6",x"44",x"58",x"CB",x"05", -- 0x8B60
    x"4F",x"33",x"CB",x"11",x"A3",x"E4",x"27",x"E2", -- 0x8B68
    x"8D",x"04",x"33",x"45",x"20",x"F5",x"AE",x"42", -- 0x8B70
    x"BC",x"09",x"48",x"24",x"0E",x"AC",x"22",x"25", -- 0x8B78
    x"0A",x"AC",x"24",x"25",x"07",x"1F",x"10",x"A3", -- 0x8B80
    x"A4",x"ED",x"42",x"39",x"6F",x"C4",x"6F",x"42", -- 0x8B88
    x"6F",x"43",x"39",x"F6",x"09",x"5B",x"5C",x"34", -- 0x8B90
    x"04",x"BD",x"C7",x"49",x"A6",x"00",x"81",x"40", -- 0x8B98
    x"26",x"0B",x"EC",x"0B",x"10",x"A3",x"24",x"25", -- 0x8BA0
    x"04",x"A3",x"A4",x"ED",x"0B",x"35",x"04",x"5A", -- 0x8BA8
    x"26",x"E5",x"35",x"56",x"11",x"B3",x"09",x"48", -- 0x8BB0
    x"27",x"06",x"A6",x"C0",x"A7",x"80",x"20",x"F4", -- 0x8BB8
    x"BF",x"09",x"48",x"BD",x"C7",x"55",x"6A",x"00", -- 0x8BC0
    x"6D",x"01",x"27",x"03",x"BD",x"C7",x"1E",x"9E", -- 0x8BC8
    x"F1",x"35",x"02",x"81",x"20",x"27",x"08",x"81", -- 0x8BD0
    x"40",x"26",x"B0",x"A6",x"0F",x"27",x"0A",x"BD", -- 0x8BD8
    x"C7",x"63",x"33",x"88",x"19",x"DF",x"EE",x"8D", -- 0x8BE0
    x"2C",x"A6",x"88",x"13",x"2A",x"9D",x"E6",x"88", -- 0x8BE8
    x"12",x"C4",x"07",x"86",x"20",x"3D",x"CE",x"06", -- 0x8BF0
    x"00",x"DF",x"EE",x"31",x"CB",x"E6",x"88",x"12", -- 0x8BF8
    x"54",x"54",x"54",x"CB",x"03",x"D7",x"ED",x"CC", -- 0x8C00
    x"11",x"02",x"97",x"EC",x"8D",x"09",x"EC",x"88", -- 0x8C08
    x"13",x"84",x"7F",x"ED",x"2E",x"C6",x"03",x"D7", -- 0x8C10
    x"EA",x"7E",x"D6",x"F2",x"0D",x"6F",x"10",x"2F", -- 0x8C18
    x"B6",x"51",x"32",x"62",x"34",x"16",x"8E",x"09", -- 0x8C20
    x"26",x"D6",x"6F",x"58",x"AE",x"85",x"E6",x"84", -- 0x8C28
    x"C1",x"10",x"27",x"36",x"81",x"0D",x"26",x"02", -- 0x8C30
    x"6F",x"06",x"81",x"20",x"25",x"02",x"6C",x"06", -- 0x8C38
    x"C1",x"40",x"26",x"1A",x"EC",x"88",x"17",x"C3", -- 0x8C40
    x"00",x"01",x"10",x"A3",x"09",x"10",x"22",x"01", -- 0x8C48
    x"7A",x"ED",x"88",x"17",x"AE",x"0B",x"30",x"8B", -- 0x8C50
    x"35",x"02",x"A7",x"1F",x"35",x"94",x"6C",x"88", -- 0x8C58
    x"18",x"E6",x"88",x"18",x"27",x"06",x"3A",x"A7", -- 0x8C60
    x"88",x"18",x"35",x"96",x"34",x"60",x"A7",x"89", -- 0x8C68
    x"01",x"18",x"E6",x"01",x"D7",x"EB",x"6C",x"04", -- 0x8C70
    x"BD",x"CB",x"DF",x"31",x"84",x"E6",x"03",x"BD", -- 0x8C78
    x"C7",x"55",x"3A",x"33",x"06",x"A6",x"24",x"81", -- 0x8C80
    x"09",x"25",x"0E",x"6A",x"24",x"6C",x"25",x"BD", -- 0x8C88
    x"C7",x"BF",x"6F",x"24",x"6F",x"25",x"A7",x"23", -- 0x8C90
    x"8C",x"8A",x"C0",x"A7",x"C4",x"30",x"A4",x"BD", -- 0x8C98
    x"C6",x"85",x"BD",x"C5",x"A9",x"35",x"60",x"35", -- 0x8CA0
    x"96",x"BD",x"D2",x"4F",x"BD",x"C7",x"9D",x"BD", -- 0x8CA8
    x"B9",x"58",x"CC",x"11",x"02",x"97",x"EC",x"D7", -- 0x8CB0
    x"EA",x"C6",x"03",x"D7",x"ED",x"8E",x"06",x"00", -- 0x8CB8
    x"9F",x"EE",x"BD",x"D6",x"F2",x"35",x"40",x"BD", -- 0x8CC0
    x"A5",x"49",x"34",x"40",x"A6",x"84",x"27",x"38", -- 0x8CC8
    x"43",x"27",x"44",x"34",x"10",x"C6",x"08",x"BD", -- 0x8CD0
    x"B9",x"A2",x"8D",x"3F",x"C6",x"03",x"BD",x"B9", -- 0x8CD8
    x"A2",x"8D",x"38",x"E6",x"00",x"C1",x"0A",x"24", -- 0x8CE0
    x"02",x"8D",x"30",x"4F",x"BD",x"BD",x"CC",x"8D", -- 0x8CE8
    x"2A",x"AE",x"E4",x"86",x"42",x"AB",x"0C",x"8D", -- 0x8CF0
    x"1F",x"E6",x"0D",x"8D",x"21",x"1F",x"89",x"4F", -- 0x8CF8
    x"BD",x"BD",x"CC",x"BD",x"B9",x"58",x"35",x"10", -- 0x8D00
    x"30",x"88",x"20",x"8C",x"07",x"00",x"25",x"B5", -- 0x8D08
    x"D6",x"ED",x"5C",x"C1",x"12",x"23",x"A4",x"39", -- 0x8D10
    x"BD",x"A2",x"82",x"7E",x"B9",x"AC",x"BD",x"C7", -- 0x8D18
    x"55",x"33",x"06",x"4F",x"4C",x"81",x"44",x"10", -- 0x8D20
    x"22",x"F9",x"28",x"30",x"C4",x"3A",x"E6",x"84", -- 0x8D28
    x"C1",x"C0",x"25",x"F0",x"39",x"0D",x"6F",x"2F", -- 0x8D30
    x"5E",x"8E",x"B0",x"69",x"AF",x"E4",x"8E",x"02", -- 0x8D38
    x"DD",x"C6",x"2C",x"D7",x"01",x"96",x"06",x"26", -- 0x8D40
    x"02",x"C6",x"20",x"8D",x"6F",x"81",x"20",x"27", -- 0x8D48
    x"FA",x"81",x"22",x"26",x"0A",x"C1",x"2C",x"26", -- 0x8D50
    x"06",x"1F",x"89",x"D7",x"01",x"20",x"22",x"C1", -- 0x8D58
    x"22",x"27",x"11",x"81",x"0D",x"26",x"0D",x"8C", -- 0x8D60
    x"02",x"DD",x"27",x"44",x"A6",x"1F",x"81",x"0A", -- 0x8D68
    x"26",x"3E",x"86",x"0D",x"4D",x"27",x"17",x"91", -- 0x8D70
    x"01",x"27",x"1D",x"34",x"04",x"A1",x"E0",x"27", -- 0x8D78
    x"17",x"A7",x"80",x"8C",x"03",x"D6",x"26",x"06", -- 0x8D80
    x"8D",x"46",x"26",x"06",x"20",x"1E",x"8D",x"40", -- 0x8D88
    x"27",x"CD",x"6F",x"84",x"8E",x"02",x"DC",x"39", -- 0x8D90
    x"81",x"22",x"27",x"04",x"81",x"20",x"26",x"F2", -- 0x8D98
    x"8D",x"2E",x"26",x"EE",x"81",x"20",x"27",x"F8", -- 0x8DA0
    x"81",x"2C",x"27",x"E6",x"81",x"0D",x"26",x"08", -- 0x8DA8
    x"8D",x"1E",x"26",x"DE",x"81",x"0A",x"27",x"DA", -- 0x8DB0
    x"8D",x"1C",x"20",x"D6",x"8D",x"12",x"27",x"15", -- 0x8DB8
    x"BD",x"C7",x"44",x"E6",x"00",x"C1",x"40",x"10", -- 0x8DC0
    x"26",x"F5",x"87",x"C6",x"4A",x"7E",x"AC",x"46", -- 0x8DC8
    x"BD",x"A1",x"76",x"0D",x"70",x"39",x"34",x"14", -- 0x8DD0
    x"BD",x"C7",x"44",x"E6",x"00",x"C1",x"40",x"26", -- 0x8DD8
    x"0B",x"EC",x"88",x"15",x"83",x"00",x"01",x"ED", -- 0x8DE0
    x"88",x"15",x"35",x"94",x"A7",x"88",x"11",x"63", -- 0x8DE8
    x"88",x"10",x"35",x"94",x"BD",x"B6",x"54",x"C1", -- 0x8DF0
    x"05",x"10",x"25",x"E6",x"4D",x"0F",x"06",x"7E", -- 0x8DF8
    x"BC",x"14",x"BD",x"B1",x"43",x"C6",x"05",x"BD", -- 0x8E00
    x"B5",x"0F",x"BD",x"BC",x"35",x"7E",x"B6",x"9B", -- 0x8E08
    x"8D",x"07",x"EC",x"07",x"DD",x"52",x"7E",x"88", -- 0x8E10
    x"0E",x"96",x"6F",x"34",x"02",x"BD",x"B1",x"43", -- 0x8E18
    x"BD",x"A5",x"AE",x"0D",x"6F",x"10",x"2F",x"E6", -- 0x8E20
    x"21",x"BD",x"C7",x"44",x"35",x"02",x"97",x"6F", -- 0x8E28
    x"6D",x"00",x"10",x"27",x"D5",x"C5",x"39",x"8D", -- 0x8E30
    x"E0",x"A6",x"01",x"97",x"EB",x"E6",x"02",x"34", -- 0x8E38
    x"10",x"BD",x"CD",x"1E",x"4A",x"C4",x"3F",x"34", -- 0x8E40
    x"04",x"1F",x"89",x"4F",x"BD",x"C7",x"79",x"EB", -- 0x8E48
    x"E0",x"89",x"00",x"35",x"10",x"34",x"02",x"A6", -- 0x8E50
    x"00",x"81",x"40",x"35",x"02",x"26",x"B5",x"34", -- 0x8E58
    x"10",x"93",x"8A",x"27",x"03",x"83",x"00",x"01", -- 0x8E60
    x"8D",x"AA",x"D6",x"4F",x"27",x"04",x"CB",x"08", -- 0x8E68
    x"D7",x"4F",x"BD",x"BC",x"5F",x"AE",x"E4",x"EC", -- 0x8E70
    x"88",x"13",x"84",x"7F",x"8D",x"96",x"0F",x"62", -- 0x8E78
    x"96",x"5C",x"D6",x"4F",x"BD",x"B9",x"C5",x"BD", -- 0x8E80
    x"BC",x"5F",x"35",x"10",x"EC",x"09",x"8D",x"84", -- 0x8E88
    x"0F",x"62",x"96",x"5C",x"D6",x"4F",x"BD",x"BB", -- 0x8E90
    x"91",x"7E",x"BC",x"EE",x"BD",x"B1",x"43",x"BD", -- 0x8E98
    x"B7",x"0E",x"C1",x"03",x"10",x"22",x"D7",x"77", -- 0x8EA0
    x"D7",x"EB",x"BD",x"C7",x"9D",x"BD",x"C7",x"55", -- 0x8EA8
    x"30",x"06",x"6F",x"E2",x"C6",x"44",x"A6",x"80", -- 0x8EB0
    x"43",x"26",x"02",x"6C",x"E4",x"5A",x"26",x"F6", -- 0x8EB8
    x"35",x"04",x"7E",x"B4",x"F3",x"BD",x"B7",x"0B", -- 0x8EC0
    x"C1",x"03",x"10",x"22",x"D7",x"51",x"F7",x"09", -- 0x8EC8
    x"5A",x"39",x"A6",x"64",x"26",x"13",x"AE",x"65", -- 0x8ED0
    x"8C",x"AF",x"9A",x"26",x"0C",x"AE",x"62",x"8C", -- 0x8ED8
    x"B1",x"66",x"26",x"05",x"8E",x"CE",x"EC",x"AF", -- 0x8EE0
    x"65",x"7E",x"88",x"46",x"35",x"02",x"46",x"BD", -- 0x8EE8
    x"B1",x"48",x"10",x"27",x"ED",x"3D",x"9E",x"52", -- 0x8EF0
    x"EC",x"02",x"10",x"83",x"09",x"89",x"25",x"07", -- 0x8EF8
    x"B3",x"09",x"4A",x"10",x"25",x"E0",x"AA",x"7E", -- 0x8F00
    x"AF",x"A4",x"81",x"CA",x"27",x"1C",x"81",x"C8", -- 0x8F08
    x"10",x"26",x"B2",x"28",x"9D",x"9F",x"81",x"2C", -- 0x8F10
    x"10",x"27",x"C7",x"34",x"BD",x"B7",x"0B",x"C1", -- 0x8F18
    x"04",x"10",x"22",x"E5",x"25",x"96",x"BC",x"7E", -- 0x8F20
    x"96",x"2E",x"BD",x"A4",x"29",x"9D",x"9F",x"7E", -- 0x8F28
    x"8C",x"1B",x"C1",x"34",x"10",x"26",x"B2",x"30", -- 0x8F30
    x"BD",x"B2",x"62",x"96",x"6F",x"34",x"02",x"BD", -- 0x8F38
    x"A5",x"AE",x"BD",x"A4",x"06",x"0D",x"6F",x"2F", -- 0x8F40
    x"13",x"BD",x"C7",x"44",x"E6",x"00",x"C1",x"40", -- 0x8F48
    x"26",x"0A",x"35",x"02",x"97",x"6F",x"EC",x"88", -- 0x8F50
    x"17",x"7E",x"B4",x"F4",x"BD",x"A3",x"5F",x"35", -- 0x8F58
    x"02",x"97",x"6F",x"D6",x"6C",x"7E",x"B4",x"F3", -- 0x8F60
    x"9D",x"9F",x"8D",x"4F",x"BD",x"83",x"6C",x"BD", -- 0x8F68
    x"83",x"6C",x"AC",x"62",x"10",x"25",x"E4",x"D2", -- 0x8F70
    x"BD",x"83",x"6C",x"BD",x"A5",x"C7",x"CC",x"02", -- 0x8F78
    x"00",x"FD",x"09",x"57",x"BD",x"CA",x"04",x"4F", -- 0x8F80
    x"8D",x"2B",x"EC",x"62",x"A3",x"64",x"C3",x"00", -- 0x8F88
    x"01",x"1F",x"02",x"8D",x"1E",x"EC",x"64",x"8D", -- 0x8F90
    x"1A",x"AE",x"64",x"A6",x"80",x"BD",x"CC",x"24", -- 0x8F98
    x"31",x"3F",x"26",x"F7",x"86",x"FF",x"8D",x"0D", -- 0x8FA0
    x"4F",x"5F",x"8D",x"07",x"35",x"36",x"8D",x"03", -- 0x8FA8
    x"7E",x"A4",x"2D",x"8D",x"00",x"BD",x"CC",x"24", -- 0x8FB0
    x"1E",x"89",x"39",x"8E",x"C2",x"AF",x"7E",x"C9", -- 0x8FB8
    x"38",x"9D",x"9F",x"8D",x"F6",x"BD",x"CA",x"07", -- 0x8FC0
    x"FC",x"09",x"57",x"83",x"02",x"00",x"10",x"26", -- 0x8FC8
    x"D6",x"44",x"9E",x"8A",x"9D",x"A5",x"27",x"06", -- 0x8FD0
    x"BD",x"B2",x"6D",x"BD",x"B7",x"3D",x"9F",x"D3", -- 0x8FD8
    x"BD",x"A5",x"C7",x"BD",x"CD",x"BC",x"34",x"02", -- 0x8FE0
    x"8D",x"29",x"1F",x"02",x"8D",x"25",x"D3",x"D3", -- 0x8FE8
    x"DD",x"9D",x"1F",x"01",x"A6",x"E0",x"10",x"26", -- 0x8FF0
    x"D4",x"33",x"BD",x"C5",x"C4",x"D6",x"70",x"27", -- 0x8FF8
    x"03",x"7E",x"C3",x"52",x"A7",x"84",x"A1",x"80", -- 0x9000
    x"27",x"03",x"7E",x"D7",x"09",x"31",x"3F",x"26", -- 0x9008
    x"E9",x"20",x"D0",x"8D",x"00",x"BD",x"CD",x"BC", -- 0x9010
    x"1E",x"89",x"39",x"9E",x"A6",x"34",x"10",x"8D", -- 0x9018
    x"35",x"96",x"EB",x"34",x"02",x"8D",x"2A",x"35", -- 0x9020
    x"02",x"91",x"EB",x"10",x"26",x"E4",x"1B",x"8D", -- 0x9028
    x"28",x"35",x"10",x"9F",x"A6",x"8D",x"1F",x"BD", -- 0x9030
    x"C6",x"8C",x"BD",x"C6",x"E5",x"8D",x"12",x"8E", -- 0x9038
    x"09",x"4C",x"FE",x"09",x"74",x"C6",x"0B",x"BD", -- 0x9040
    x"A5",x"9A",x"C6",x"03",x"D7",x"EA",x"7E",x"D6", -- 0x9048
    x"F2",x"C6",x"A5",x"BD",x"B2",x"6F",x"7E",x"C9", -- 0x9050
    x"35",x"BD",x"C6",x"8C",x"C6",x"42",x"7D",x"09", -- 0x9058
    x"73",x"10",x"26",x"DB",x"E1",x"39",x"10",x"27", -- 0x9060
    x"E8",x"EE",x"8D",x"03",x"0F",x"6F",x"39",x"81", -- 0x9068
    x"23",x"26",x"0F",x"BD",x"A5",x"A5",x"BD",x"A4", -- 0x9070
    x"06",x"9D",x"A5",x"10",x"27",x"E8",x"D9",x"BD", -- 0x9078
    x"B2",x"6D",x"BD",x"B1",x"56",x"96",x"06",x"26", -- 0x9080
    x"1E",x"BD",x"BD",x"D9",x"BD",x"B5",x"16",x"BD", -- 0x9088
    x"B9",x"9F",x"9D",x"A5",x"10",x"27",x"E8",x"C0", -- 0x9090
    x"86",x"2C",x"BD",x"A3",x"5F",x"0D",x"6E",x"27", -- 0x9098
    x"02",x"86",x"0D",x"8D",x"14",x"20",x"D8",x"8D", -- 0x90A0
    x"07",x"BD",x"B9",x"9F",x"8D",x"02",x"20",x"E2", -- 0x90A8
    x"BD",x"A3",x"5F",x"0D",x"6E",x"26",x"B7",x"86", -- 0x90B0
    x"22",x"7E",x"A2",x"82",x"BD",x"C8",x"2E",x"4F", -- 0x90B8
    x"5F",x"34",x"16",x"9D",x"A5",x"26",x"02",x"35", -- 0x90C0
    x"96",x"BD",x"B7",x"38",x"34",x"14",x"4F",x"E3", -- 0x90C8
    x"63",x"25",x"07",x"AE",x"65",x"10",x"A3",x"09", -- 0x90D0
    x"23",x"05",x"C6",x"44",x"7E",x"AC",x"46",x"EE", -- 0x90D8
    x"63",x"ED",x"63",x"EC",x"0B",x"33",x"CB",x"EF", -- 0x90E0
    x"61",x"C6",x"FF",x"BD",x"B2",x"6F",x"C6",x"A7", -- 0x90E8
    x"BD",x"B2",x"6F",x"BD",x"B3",x"57",x"BD",x"B1", -- 0x90F0
    x"46",x"35",x"44",x"E7",x"84",x"EF",x"02",x"20", -- 0x90F8
    x"C2",x"86",x"4F",x"34",x"02",x"BD",x"B3",x"57", -- 0x9100
    x"BD",x"B1",x"46",x"34",x"10",x"AE",x"02",x"8C", -- 0x9108
    x"09",x"89",x"25",x"05",x"BC",x"09",x"4A",x"25", -- 0x9110
    x"05",x"C6",x"46",x"7E",x"AC",x"46",x"C6",x"B3", -- 0x9118
    x"BD",x"B2",x"6F",x"BD",x"87",x"48",x"35",x"20", -- 0x9120
    x"A6",x"A4",x"27",x"2E",x"34",x"04",x"C6",x"20", -- 0x9128
    x"EE",x"22",x"E7",x"C0",x"4A",x"26",x"FB",x"E6", -- 0x9130
    x"E0",x"27",x"1F",x"E1",x"A4",x"25",x"04",x"E6", -- 0x9138
    x"A4",x"6F",x"E4",x"EE",x"22",x"6D",x"E0",x"27", -- 0x9140
    x"0E",x"34",x"04",x"4F",x"50",x"82",x"00",x"EB", -- 0x9148
    x"A4",x"89",x"00",x"33",x"CB",x"35",x"04",x"7E", -- 0x9150
    x"A5",x"9A",x"35",x"82",x"BD",x"95",x"AC",x"FC", -- 0x9158
    x"09",x"4A",x"83",x"09",x"89",x"34",x"06",x"F6", -- 0x9160
    x"09",x"5B",x"34",x"04",x"9D",x"A5",x"81",x"2C", -- 0x9168
    x"27",x"0F",x"BD",x"B7",x"0B",x"C1",x"0F",x"10", -- 0x9170
    x"22",x"E2",x"CF",x"E7",x"E4",x"9D",x"A5",x"27", -- 0x9178
    x"08",x"BD",x"B2",x"6D",x"BD",x"B3",x"E6",x"ED", -- 0x9180
    x"61",x"BD",x"CA",x"E9",x"E6",x"E4",x"34",x"04", -- 0x9188
    x"CC",x"09",x"89",x"E3",x"62",x"25",x"71",x"ED", -- 0x9190
    x"62",x"C3",x"01",x"19",x"25",x"6A",x"6A",x"E4", -- 0x9198
    x"2A",x"F7",x"5D",x"27",x"03",x"4C",x"27",x"60", -- 0x91A0
    x"85",x"01",x"27",x"03",x"4C",x"27",x"59",x"A7", -- 0x91A8
    x"E4",x"DC",x"1B",x"90",x"BC",x"AB",x"E4",x"25", -- 0x91B0
    x"4F",x"1F",x"01",x"4C",x"27",x"4A",x"10",x"93", -- 0x91B8
    x"21",x"24",x"45",x"4A",x"93",x"1B",x"D3",x"19", -- 0x91C0
    x"1F",x"02",x"A6",x"E4",x"90",x"BC",x"1F",x"89", -- 0x91C8
    x"9B",x"BA",x"97",x"BA",x"DB",x"B7",x"D7",x"B7", -- 0x91D0
    x"35",x"46",x"97",x"BC",x"F7",x"09",x"5B",x"FF", -- 0x91D8
    x"09",x"4A",x"96",x"68",x"4C",x"27",x"08",x"1F", -- 0x91E0
    x"20",x"93",x"19",x"D3",x"A6",x"DD",x"A6",x"DE", -- 0x91E8
    x"1B",x"9F",x"1B",x"11",x"93",x"1B",x"22",x"13", -- 0x91F0
    x"A6",x"C2",x"A7",x"82",x"11",x"93",x"19",x"26", -- 0x91F8
    x"F7",x"10",x"9F",x"19",x"6F",x"3F",x"20",x"13", -- 0x9200
    x"7E",x"AC",x"44",x"DE",x"19",x"10",x"9F",x"19", -- 0x9208
    x"6F",x"3F",x"A6",x"C0",x"A7",x"A0",x"10",x"9C", -- 0x9210
    x"1B",x"26",x"F7",x"CE",x"09",x"28",x"BE",x"09", -- 0x9218
    x"4A",x"5F",x"AF",x"C1",x"6F",x"00",x"30",x"89", -- 0x9220
    x"01",x"19",x"5C",x"F1",x"09",x"5B",x"23",x"F2", -- 0x9228
    x"7E",x"96",x"CB",x"8D",x"1A",x"5F",x"5C",x"BD", -- 0x9230
    x"C7",x"49",x"27",x"0D",x"A6",x"01",x"91",x"EB", -- 0x9238
    x"26",x"07",x"34",x"04",x"BD",x"CB",x"06",x"35", -- 0x9240
    x"04",x"F1",x"09",x"5B",x"23",x"E8",x"39",x"F6", -- 0x9248
    x"09",x"5A",x"9D",x"A5",x"27",x"09",x"BD",x"B7", -- 0x9250
    x"0B",x"C1",x"03",x"10",x"22",x"D3",x"C0",x"D7", -- 0x9258
    x"EB",x"39",x"10",x"27",x"D3",x"B9",x"BD",x"95", -- 0x9260
    x"AC",x"BD",x"D2",x"56",x"F7",x"06",x"FF",x"9D", -- 0x9268
    x"A5",x"27",x"08",x"C6",x"A5",x"BD",x"B2",x"6F", -- 0x9270
    x"BD",x"D2",x"56",x"10",x"CE",x"06",x"FF",x"34", -- 0x9278
    x"04",x"BD",x"A5",x"C7",x"BD",x"CA",x"E9",x"6F", -- 0x9280
    x"E2",x"8E",x"09",x"88",x"6C",x"E4",x"30",x"89", -- 0x9288
    x"12",x"00",x"9C",x"27",x"23",x"F6",x"6A",x"E4", -- 0x9290
    x"10",x"27",x"D9",x"A8",x"86",x"23",x"5F",x"34", -- 0x9298
    x"06",x"73",x"09",x"5C",x"5F",x"5C",x"6A",x"E4", -- 0x92A0
    x"27",x"04",x"E1",x"62",x"26",x"F7",x"D7",x"03", -- 0x92A8
    x"E6",x"64",x"8D",x"48",x"86",x"FF",x"BD",x"D3", -- 0x92B0
    x"22",x"E6",x"63",x"8D",x"42",x"6D",x"E4",x"27", -- 0x92B8
    x"0C",x"4F",x"BD",x"D3",x"22",x"E6",x"61",x"DB", -- 0x92C0
    x"03",x"E7",x"61",x"20",x"D7",x"8D",x"03",x"7E", -- 0x92C8
    x"AC",x"73",x"35",x"40",x"B6",x"09",x"5C",x"27", -- 0x92D0
    x"16",x"8E",x"09",x"28",x"4F",x"6F",x"91",x"4C", -- 0x92D8
    x"B1",x"09",x"5B",x"23",x"F8",x"9E",x"19",x"6F", -- 0x92E0
    x"1F",x"BD",x"AD",x"19",x"7F",x"09",x"5C",x"B6", -- 0x92E8
    x"09",x"5D",x"27",x"06",x"7F",x"09",x"5D",x"BD", -- 0x92F0
    x"AD",x"19",x"6E",x"C4",x"86",x"02",x"8C",x"86", -- 0x92F8
    x"03",x"DD",x"EA",x"A6",x"63",x"97",x"EC",x"8E", -- 0x9300
    x"09",x"89",x"9F",x"EE",x"96",x"03",x"C6",x"01", -- 0x9308
    x"D7",x"ED",x"BD",x"D6",x"F2",x"0C",x"EE",x"5C", -- 0x9310
    x"C1",x"12",x"23",x"F4",x"0C",x"EC",x"4A",x"26", -- 0x9318
    x"ED",x"39",x"E6",x"65",x"E1",x"66",x"26",x"36", -- 0x9320
    x"7F",x"09",x"85",x"7F",x"FF",x"40",x"7F",x"09", -- 0x9328
    x"86",x"34",x"02",x"BD",x"A9",x"28",x"8E",x"D3", -- 0x9330
    x"5F",x"C6",x"0D",x"A6",x"E0",x"27",x"05",x"8E", -- 0x9338
    x"D3",x"6C",x"C6",x"12",x"BD",x"B9",x"A2",x"8E", -- 0x9340
    x"D3",x"7E",x"C6",x"1B",x"BD",x"B9",x"A2",x"CC", -- 0x9348
    x"64",x"05",x"97",x"8C",x"BD",x"A9",x"51",x"BD", -- 0x9350
    x"A1",x"71",x"81",x"0D",x"26",x"F9",x"39",x"49", -- 0x9358
    x"4E",x"53",x"45",x"52",x"54",x"20",x"53",x"4F", -- 0x9360
    x"55",x"52",x"43",x"45",x"49",x"4E",x"53",x"45", -- 0x9368
    x"52",x"54",x"20",x"44",x"45",x"53",x"54",x"49", -- 0x9370
    x"4E",x"41",x"54",x"49",x"4F",x"4E",x"20",x"44", -- 0x9378
    x"49",x"53",x"4B",x"45",x"54",x"54",x"45",x"20", -- 0x9380
    x"41",x"4E",x"44",x"0D",x"50",x"52",x"45",x"53", -- 0x9388
    x"53",x"20",x"27",x"45",x"4E",x"54",x"45",x"52", -- 0x9390
    x"27",x"35",x"20",x"C6",x"0B",x"8E",x"09",x"57", -- 0x9398
    x"A6",x"82",x"34",x"02",x"5A",x"26",x"F9",x"96", -- 0x93A0
    x"EB",x"34",x"02",x"6E",x"A4",x"A6",x"80",x"97", -- 0x93A8
    x"EB",x"C6",x"0B",x"CE",x"09",x"4C",x"7E",x"A5", -- 0x93B0
    x"9A",x"BD",x"C9",x"35",x"8D",x"DB",x"6F",x"E2", -- 0x93B8
    x"9D",x"A5",x"27",x"0A",x"63",x"E4",x"C6",x"A5", -- 0x93C0
    x"BD",x"B2",x"6F",x"BD",x"C9",x"35",x"8D",x"C9", -- 0x93C8
    x"BD",x"A5",x"C7",x"BD",x"CA",x"E9",x"6F",x"E2", -- 0x93D0
    x"30",x"E9",x"FF",x"00",x"6C",x"E4",x"30",x"89", -- 0x93D8
    x"FF",x"00",x"9C",x"1F",x"24",x"F6",x"6A",x"E4", -- 0x93E0
    x"10",x"27",x"D8",x"58",x"30",x"6E",x"8D",x"BD", -- 0x93E8
    x"BD",x"C6",x"8C",x"BD",x"C6",x"E5",x"BE",x"09", -- 0x93F0
    x"74",x"EE",x"0E",x"AE",x"0B",x"34",x"50",x"BD", -- 0x93F8
    x"C7",x"9D",x"F6",x"09",x"76",x"BD",x"CD",x"1E", -- 0x9400
    x"34",x"02",x"4A",x"C4",x"3F",x"34",x"04",x"1F", -- 0x9408
    x"89",x"4F",x"BD",x"C7",x"79",x"EB",x"E4",x"89", -- 0x9410
    x"00",x"8E",x"00",x"01",x"34",x"16",x"5F",x"AE", -- 0x9418
    x"E4",x"27",x"09",x"5C",x"30",x"1F",x"27",x"04", -- 0x9420
    x"E1",x"6A",x"26",x"F7",x"AF",x"E4",x"E7",x"64", -- 0x9428
    x"8D",x"50",x"86",x"FF",x"8D",x"40",x"6D",x"65", -- 0x9430
    x"27",x"25",x"30",x"6B",x"BD",x"D3",x"AD",x"BD", -- 0x9438
    x"D0",x"59",x"BD",x"C7",x"9D",x"BD",x"C7",x"55", -- 0x9440
    x"30",x"06",x"A6",x"65",x"C6",x"44",x"63",x"84", -- 0x9448
    x"26",x"03",x"4A",x"27",x"08",x"63",x"80",x"5A", -- 0x9450
    x"26",x"F4",x"7E",x"C7",x"F8",x"63",x"84",x"8D", -- 0x9458
    x"1B",x"AE",x"E4",x"27",x"0D",x"EC",x"62",x"EB", -- 0x9460
    x"64",x"89",x"00",x"ED",x"62",x"4F",x"8D",x"06", -- 0x9468
    x"20",x"AC",x"32",x"E8",x"24",x"39",x"6D",x"E8", -- 0x9470
    x"19",x"7E",x"D3",x"26",x"86",x"FF",x"30",x"6D", -- 0x9478
    x"20",x"04",x"4F",x"30",x"E8",x"1A",x"97",x"D8", -- 0x9480
    x"BD",x"D3",x"AD",x"AE",x"68",x"BF",x"09",x"57", -- 0x9488
    x"8E",x"01",x"00",x"BF",x"09",x"7C",x"86",x"52", -- 0x9490
    x"F6",x"09",x"5B",x"5C",x"BD",x"C4",x"8D",x"9E", -- 0x9498
    x"F1",x"CC",x"01",x"00",x"ED",x"88",x"13",x"E6", -- 0x94A0
    x"66",x"27",x"29",x"D6",x"D8",x"E4",x"67",x"27", -- 0x94A8
    x"09",x"EC",x"62",x"EB",x"66",x"89",x"00",x"BD", -- 0x94B0
    x"C2",x"E6",x"9E",x"F1",x"EE",x"64",x"EF",x"07", -- 0x94B8
    x"E6",x"66",x"DE",x"1F",x"34",x"44",x"9E",x"F1", -- 0x94C0
    x"EF",x"0B",x"BD",x"C2",x"EA",x"6C",x"61",x"35", -- 0x94C8
    x"44",x"5A",x"26",x"F0",x"9E",x"F1",x"CE",x"09", -- 0x94D0
    x"89",x"EF",x"0B",x"D6",x"D8",x"E4",x"67",x"27", -- 0x94D8
    x"09",x"6F",x"67",x"EC",x"6A",x"8A",x"80",x"ED", -- 0x94E0
    x"88",x"13",x"7E",x"CB",x"06",x"8D",x"38",x"8D", -- 0x94E8
    x"2B",x"34",x"10",x"8D",x"27",x"34",x"10",x"C6", -- 0x94F0
    x"02",x"BD",x"D5",x"8F",x"CE",x"06",x"80",x"35", -- 0x94F8
    x"10",x"8D",x"05",x"CE",x"06",x"00",x"35",x"10", -- 0x9500
    x"34",x"50",x"C6",x"80",x"BD",x"B5",x"0F",x"33", -- 0x9508
    x"84",x"35",x"10",x"E7",x"84",x"EF",x"02",x"35", -- 0x9510
    x"10",x"7E",x"A5",x"9A",x"BD",x"B2",x"6D",x"8E", -- 0x9518
    x"B3",x"57",x"8D",x"2F",x"7E",x"B1",x"46",x"BD", -- 0x9520
    x"B7",x"0B",x"C1",x"03",x"22",x"1C",x"34",x"04", -- 0x9528
    x"BD",x"B7",x"38",x"C1",x"22",x"22",x"13",x"34", -- 0x9530
    x"04",x"BD",x"B7",x"38",x"D7",x"ED",x"5A",x"C1", -- 0x9538
    x"11",x"22",x"07",x"35",x"06",x"97",x"EC",x"D7", -- 0x9540
    x"EB",x"39",x"7E",x"B4",x"4A",x"BD",x"B2",x"6D", -- 0x9548
    x"8E",x"B1",x"56",x"D6",x"EB",x"DE",x"EC",x"34", -- 0x9550
    x"44",x"AD",x"84",x"35",x"44",x"D7",x"EB",x"DF", -- 0x9558
    x"EC",x"39",x"8D",x"C3",x"8D",x"E7",x"8D",x"BC", -- 0x9560
    x"9E",x"52",x"34",x"10",x"8D",x"DF",x"BD",x"B6", -- 0x9568
    x"54",x"34",x"14",x"5F",x"8E",x"06",x"00",x"6F", -- 0x9570
    x"80",x"5A",x"26",x"FB",x"35",x"14",x"CE",x"06", -- 0x9578
    x"80",x"8D",x"96",x"35",x"10",x"BD",x"B6",x"59", -- 0x9580
    x"CE",x"06",x"00",x"8D",x"8C",x"C6",x"03",x"8E", -- 0x9588
    x"06",x"00",x"9F",x"EE",x"D7",x"EA",x"7E",x"D6", -- 0x9590
    x"F2",x"10",x"27",x"D0",x"82",x"BD",x"D2",x"56", -- 0x9598
    x"C6",x"04",x"9D",x"A5",x"27",x"0C",x"BD",x"B7", -- 0x95A0
    x"38",x"C1",x"11",x"10",x"24",x"DE",x"9B",x"BD", -- 0x95A8
    x"A5",x"C7",x"34",x"04",x"8E",x"07",x"12",x"C6", -- 0x95B0
    x"12",x"6F",x"82",x"5A",x"26",x"FB",x"4F",x"20", -- 0x95B8
    x"0D",x"EB",x"E4",x"5C",x"C0",x"12",x"24",x"FC", -- 0x95C0
    x"CB",x"12",x"6D",x"85",x"26",x"F5",x"4C",x"A7", -- 0x95C8
    x"85",x"81",x"12",x"25",x"EC",x"32",x"61",x"8E", -- 0x95D0
    x"22",x"0F",x"9C",x"27",x"10",x"22",x"D6",x"64", -- 0x95D8
    x"BD",x"CA",x"E9",x"73",x"09",x"5C",x"10",x"CE", -- 0x95E0
    x"08",x"00",x"BD",x"95",x"AC",x"86",x"00",x"97", -- 0x95E8
    x"EA",x"0F",x"EC",x"BD",x"D6",x"F2",x"7F",x"09", -- 0x95F0
    x"85",x"86",x"C0",x"B7",x"FF",x"48",x"BD",x"D7", -- 0x95F8
    x"D1",x"27",x"1D",x"7E",x"D6",x"88",x"81",x"16", -- 0x9600
    x"25",x"08",x"B6",x"09",x"86",x"8A",x"10",x"B7", -- 0x9608
    x"FF",x"40",x"86",x"53",x"B7",x"FF",x"48",x"1E", -- 0x9610
    x"88",x"1E",x"88",x"BD",x"D7",x"D1",x"26",x"68", -- 0x9618
    x"BD",x"D7",x"F0",x"8D",x"6C",x"10",x"8E",x"FF", -- 0x9620
    x"4B",x"1A",x"50",x"8E",x"D6",x"4F",x"BF",x"09", -- 0x9628
    x"83",x"8E",x"09",x"89",x"B6",x"FF",x"48",x"86", -- 0x9630
    x"FF",x"B7",x"09",x"82",x"C6",x"F4",x"F7",x"FF", -- 0x9638
    x"48",x"B6",x"09",x"86",x"8A",x"80",x"B7",x"FF", -- 0x9640
    x"40",x"E6",x"80",x"E7",x"A4",x"20",x"FA",x"B6", -- 0x9648
    x"FF",x"48",x"1C",x"AF",x"84",x"44",x"97",x"F0", -- 0x9650
    x"26",x"2E",x"0C",x"EC",x"96",x"EC",x"81",x"23", -- 0x9658
    x"26",x"A4",x"86",x"02",x"97",x"EA",x"8E",x"06", -- 0x9660
    x"00",x"9F",x"EE",x"CE",x"07",x"00",x"4F",x"97", -- 0x9668
    x"EC",x"5F",x"A6",x"C5",x"97",x"ED",x"BD",x"D6", -- 0x9670
    x"F2",x"5C",x"C1",x"12",x"25",x"F4",x"96",x"EC", -- 0x9678
    x"4C",x"81",x"23",x"25",x"EA",x"7E",x"D2",x"CD", -- 0x9680
    x"7F",x"09",x"86",x"7F",x"FF",x"40",x"7E",x"D7", -- 0x9688
    x"01",x"8E",x"09",x"89",x"CC",x"20",x"4E",x"8D", -- 0x9690
    x"29",x"5F",x"34",x"04",x"CE",x"07",x"00",x"E6", -- 0x9698
    x"C5",x"D7",x"ED",x"CE",x"D6",x"D4",x"C6",x"03", -- 0x96A0
    x"8D",x"1E",x"96",x"EC",x"A7",x"80",x"6F",x"80", -- 0x96A8
    x"96",x"ED",x"A7",x"80",x"C6",x"09",x"8D",x"10", -- 0x96B0
    x"35",x"04",x"5C",x"C1",x"12",x"25",x"DB",x"CC", -- 0x96B8
    x"C8",x"4E",x"E7",x"80",x"4A",x"26",x"FB",x"39", -- 0x96C0
    x"34",x"04",x"EC",x"C1",x"8D",x"F4",x"35",x"04", -- 0x96C8
    x"5A",x"26",x"F5",x"39",x"08",x"00",x"03",x"F5", -- 0x96D0
    x"01",x"FE",x"01",x"01",x"01",x"F7",x"16",x"4E", -- 0x96D8
    x"0C",x"00",x"03",x"F5",x"01",x"FB",x"00",x"FF", -- 0x96E0
    x"01",x"F7",x"18",x"4E",x"26",x"54",x"6E",x"9F", -- 0x96E8
    x"C0",x"0A",x"34",x"04",x"C6",x"05",x"F7",x"09", -- 0x96F0
    x"88",x"35",x"04",x"8D",x"62",x"0D",x"F0",x"27", -- 0x96F8
    x"0D",x"96",x"F0",x"C6",x"3C",x"85",x"40",x"26", -- 0x9700
    x"02",x"C6",x"28",x"7E",x"AC",x"46",x"34",x"02", -- 0x9708
    x"96",x"EA",x"81",x"03",x"35",x"02",x"26",x"2A", -- 0x9710
    x"7D",x"09",x"87",x"27",x"25",x"34",x"56",x"86", -- 0x9718
    x"02",x"97",x"EA",x"DE",x"EE",x"8E",x"07",x"00", -- 0x9720
    x"9F",x"EE",x"8D",x"33",x"DF",x"EE",x"86",x"03", -- 0x9728
    x"97",x"EA",x"96",x"F0",x"26",x"0D",x"5F",x"A6", -- 0x9730
    x"80",x"A1",x"C0",x"26",x"06",x"5A",x"26",x"F7", -- 0x9738
    x"35",x"56",x"39",x"35",x"56",x"7A",x"09",x"88", -- 0x9740
    x"26",x"B1",x"C6",x"48",x"20",x"BD",x"5F",x"81", -- 0x9748
    x"AA",x"27",x"07",x"53",x"81",x"88",x"10",x"26", -- 0x9750
    x"DB",x"1D",x"F7",x"09",x"87",x"0E",x"9F",x"34", -- 0x9758
    x"76",x"86",x"05",x"34",x"02",x"7F",x"09",x"85", -- 0x9760
    x"D6",x"EB",x"8E",x"D8",x"9D",x"B6",x"09",x"86", -- 0x9768
    x"84",x"A8",x"AA",x"85",x"8A",x"20",x"D6",x"EC", -- 0x9770
    x"C1",x"16",x"25",x"02",x"8A",x"10",x"1F",x"89", -- 0x9778
    x"8A",x"08",x"B7",x"09",x"86",x"B7",x"FF",x"40", -- 0x9780
    x"C5",x"08",x"26",x"06",x"BD",x"A7",x"D1",x"BD", -- 0x9788
    x"A7",x"D1",x"8D",x"3D",x"26",x"0A",x"0F",x"F0", -- 0x9790
    x"8E",x"D8",x"95",x"D6",x"EA",x"58",x"AD",x"95", -- 0x9798
    x"35",x"02",x"D6",x"F0",x"27",x"0B",x"4A",x"27", -- 0x97A0
    x"08",x"34",x"02",x"8D",x"0B",x"26",x"F1",x"20", -- 0x97A8
    x"B4",x"86",x"78",x"B7",x"09",x"85",x"35",x"F6", -- 0x97B0
    x"8E",x"09",x"7E",x"D6",x"EB",x"6F",x"85",x"86", -- 0x97B8
    x"03",x"B7",x"FF",x"48",x"1E",x"88",x"1E",x"88", -- 0x97C0
    x"8D",x"07",x"8D",x"24",x"84",x"10",x"97",x"F0", -- 0x97C8
    x"39",x"9E",x"8A",x"30",x"1F",x"27",x"08",x"B6", -- 0x97D0
    x"FF",x"48",x"85",x"01",x"26",x"F5",x"39",x"86", -- 0x97D8
    x"D0",x"B7",x"FF",x"48",x"1E",x"88",x"1E",x"88", -- 0x97E0
    x"B6",x"FF",x"48",x"86",x"80",x"97",x"F0",x"39", -- 0x97E8
    x"8E",x"22",x"2E",x"30",x"1F",x"26",x"FC",x"39", -- 0x97F0
    x"86",x"80",x"8C",x"86",x"A0",x"34",x"02",x"8E", -- 0x97F8
    x"09",x"7E",x"D6",x"EB",x"3A",x"E6",x"84",x"F7", -- 0x9800
    x"FF",x"49",x"D1",x"EC",x"27",x"1E",x"96",x"EC", -- 0x9808
    x"B7",x"FF",x"4B",x"A7",x"84",x"86",x"17",x"B7", -- 0x9810
    x"FF",x"48",x"1E",x"88",x"1E",x"88",x"8D",x"B1", -- 0x9818
    x"26",x"08",x"8D",x"CC",x"84",x"18",x"27",x"04", -- 0x9820
    x"97",x"F0",x"35",x"82",x"96",x"ED",x"B7",x"FF", -- 0x9828
    x"4A",x"8E",x"D8",x"8B",x"BF",x"09",x"83",x"9E", -- 0x9830
    x"EE",x"B6",x"FF",x"48",x"B6",x"09",x"86",x"8A", -- 0x9838
    x"80",x"35",x"04",x"10",x"9E",x"8A",x"CE",x"FF", -- 0x9840
    x"48",x"73",x"09",x"82",x"1A",x"50",x"F7",x"FF", -- 0x9848
    x"48",x"1E",x"88",x"1E",x"88",x"C1",x"80",x"27", -- 0x9850
    x"1C",x"C6",x"02",x"E5",x"C4",x"26",x"0C",x"31", -- 0x9858
    x"3F",x"26",x"F8",x"7F",x"09",x"82",x"1C",x"AF", -- 0x9860
    x"7E",x"D7",x"DF",x"E6",x"80",x"F7",x"FF",x"4B", -- 0x9868
    x"B7",x"FF",x"40",x"20",x"F6",x"C6",x"02",x"E5", -- 0x9870
    x"C4",x"26",x"06",x"31",x"3F",x"26",x"F8",x"20", -- 0x9878
    x"E2",x"F6",x"FF",x"4B",x"E7",x"80",x"B7",x"FF", -- 0x9880
    x"40",x"20",x"F6",x"1C",x"AF",x"B6",x"FF",x"48", -- 0x9888
    x"84",x"7C",x"97",x"F0",x"39",x"D7",x"B8",x"D7", -- 0x9890
    x"D0",x"D7",x"F8",x"D7",x"FB",x"01",x"02",x"04", -- 0x9898
    x"40",x"B6",x"09",x"82",x"27",x"08",x"BE",x"09", -- 0x98A0
    x"83",x"AF",x"6A",x"7F",x"09",x"82",x"3B",x"B6", -- 0x98A8
    x"FF",x"03",x"2A",x"FA",x"B6",x"FF",x"02",x"B6", -- 0x98B0
    x"09",x"85",x"27",x"11",x"4A",x"B7",x"09",x"85", -- 0x98B8
    x"26",x"0B",x"B6",x"09",x"86",x"84",x"B0",x"B7", -- 0x98C0
    x"09",x"86",x"B7",x"FF",x"40",x"7E",x"89",x"55", -- 0x98C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x98D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x98D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x98E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x98E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x98F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x98F8
    x"13",x"34",x"06",x"9D",x"A5",x"27",x"03",x"BD", -- 0x9900
    x"95",x"81",x"96",x"B5",x"97",x"D8",x"35",x"06", -- 0x9908
    x"DD",x"B4",x"4F",x"34",x"56",x"BD",x"95",x"22", -- 0x9910
    x"BD",x"92",x"8F",x"DF",x"D9",x"BD",x"99",x"DF", -- 0x9918
    x"27",x"0F",x"BD",x"99",x"CB",x"86",x"01",x"97", -- 0x9920
    x"D7",x"BD",x"99",x"BA",x"00",x"D7",x"BD",x"99", -- 0x9928
    x"BA",x"10",x"DF",x"DC",x"0D",x"DB",x"26",x"03", -- 0x9930
    x"10",x"DE",x"DC",x"35",x"56",x"0F",x"DB",x"10", -- 0x9938
    x"DF",x"DC",x"30",x"01",x"9F",x"BD",x"DF",x"D1", -- 0x9940
    x"97",x"D7",x"27",x"9F",x"2B",x"06",x"5C",x"D1", -- 0x9948
    x"D6",x"23",x"05",x"5F",x"5D",x"27",x"DD",x"5A", -- 0x9950
    x"D7",x"C0",x"BD",x"99",x"DF",x"27",x"0F",x"10", -- 0x9958
    x"83",x"00",x"03",x"25",x"04",x"30",x"1E",x"8D", -- 0x9960
    x"38",x"BD",x"99",x"CB",x"8D",x"4C",x"43",x"53", -- 0x9968
    x"D3",x"D1",x"DD",x"D1",x"2F",x"16",x"BD",x"95", -- 0x9970
    x"06",x"BD",x"9A",x"12",x"26",x"05",x"CC",x"FF", -- 0x9978
    x"FF",x"20",x"ED",x"BD",x"95",x"14",x"8D",x"3E", -- 0x9980
    x"8D",x"5E",x"20",x"E0",x"BD",x"95",x"06",x"30", -- 0x9988
    x"8B",x"9F",x"BD",x"43",x"53",x"83",x"00",x"01", -- 0x9990
    x"2F",x"04",x"1F",x"01",x"8D",x"03",x"7E",x"99", -- 0x9998
    x"34",x"DD",x"CB",x"35",x"20",x"DC",x"BD",x"34", -- 0x99A0
    x"16",x"96",x"D7",x"40",x"D6",x"C0",x"34",x"06", -- 0x99A8
    x"34",x"20",x"C6",x"02",x"BD",x"AC",x"33",x"DC", -- 0x99B0
    x"CB",x"39",x"DD",x"CB",x"35",x"20",x"DC",x"C3", -- 0x99B8
    x"34",x"16",x"96",x"D7",x"20",x"E6",x"9E",x"BD", -- 0x99C0
    x"9F",x"C3",x"39",x"DD",x"CD",x"10",x"9E",x"C3", -- 0x99C8
    x"8D",x"F4",x"10",x"9F",x"BD",x"8D",x"11",x"9E", -- 0x99D0
    x"CD",x"30",x"8B",x"C3",x"00",x"01",x"39",x"BD", -- 0x99D8
    x"99",x"C6",x"10",x"8E",x"95",x"14",x"20",x"06", -- 0x99E0
    x"10",x"8E",x"95",x"06",x"AD",x"A4",x"DE",x"8A", -- 0x99E8
    x"9E",x"BD",x"2B",x"17",x"9C",x"D3",x"22",x"13", -- 0x99F0
    x"34",x"60",x"8D",x"16",x"27",x"0B",x"BD",x"93", -- 0x99F8
    x"77",x"35",x"60",x"33",x"41",x"AD",x"A4",x"20", -- 0x9A00
    x"E9",x"35",x"60",x"1F",x"30",x"1F",x"01",x"93", -- 0x9A08
    x"8A",x"39",x"AD",x"9F",x"00",x"D9",x"1F",x"89", -- 0x9A10
    x"D4",x"D8",x"34",x"06",x"A4",x"84",x"A1",x"61", -- 0x9A18
    x"35",x"86",x"9E",x"8A",x"C6",x"01",x"34",x"14", -- 0x9A20
    x"BD",x"B1",x"56",x"5F",x"BD",x"A9",x"A2",x"BD", -- 0x9A28
    x"A9",x"76",x"BD",x"B6",x"54",x"20",x"02",x"35", -- 0x9A30
    x"14",x"D7",x"D8",x"27",x"FA",x"9F",x"D9",x"10", -- 0x9A38
    x"27",x"0F",x"31",x"0D",x"D8",x"27",x"F0",x"BD", -- 0x9A40
    x"9B",x"98",x"81",x"3B",x"27",x"F5",x"81",x"27", -- 0x9A48
    x"27",x"F1",x"81",x"58",x"10",x"27",x"01",x"B2", -- 0x9A50
    x"8D",x"02",x"20",x"E7",x"81",x"4F",x"26",x"0D", -- 0x9A58
    x"D6",x"DE",x"5C",x"8D",x"5B",x"5A",x"C1",x"04", -- 0x9A60
    x"22",x"63",x"D7",x"DE",x"39",x"81",x"56",x"26", -- 0x9A68
    x"1A",x"D6",x"DF",x"54",x"54",x"C0",x"1F",x"8D", -- 0x9A70
    x"47",x"C1",x"1F",x"22",x"50",x"58",x"58",x"34", -- 0x9A78
    x"04",x"CC",x"7E",x"7E",x"AB",x"E4",x"E0",x"E0", -- 0x9A80
    x"DD",x"DF",x"39",x"81",x"4C",x"26",x"23",x"D6", -- 0x9A88
    x"E1",x"8D",x"2D",x"5D",x"27",x"37",x"D7",x"E1", -- 0x9A90
    x"0F",x"E5",x"8D",x"03",x"24",x"FC",x"39",x"0D", -- 0x9A98
    x"D8",x"27",x"0A",x"BD",x"9B",x"98",x"81",x"2E", -- 0x9AA0
    x"27",x"05",x"BD",x"9B",x"E2",x"43",x"39",x"0C", -- 0x9AA8
    x"E5",x"39",x"81",x"54",x"26",x"0D",x"D6",x"E2", -- 0x9AB0
    x"8D",x"06",x"5D",x"27",x"10",x"D7",x"E2",x"39", -- 0x9AB8
    x"7E",x"9B",x"AC",x"81",x"50",x"26",x"24",x"BD", -- 0x9AC0
    x"9C",x"CB",x"5D",x"26",x"03",x"7E",x"B4",x"4A", -- 0x9AC8
    x"96",x"E5",x"9E",x"DF",x"34",x"12",x"86",x"7E", -- 0x9AD0
    x"97",x"DF",x"97",x"E0",x"0F",x"E5",x"8D",x"07", -- 0x9AD8
    x"35",x"12",x"97",x"E5",x"9F",x"DF",x"39",x"6F", -- 0x9AE0
    x"E2",x"20",x"40",x"81",x"4E",x"26",x"03",x"BD", -- 0x9AE8
    x"9B",x"98",x"81",x"41",x"25",x"04",x"81",x"47", -- 0x9AF0
    x"23",x"05",x"BD",x"9B",x"BE",x"20",x"23",x"80", -- 0x9AF8
    x"41",x"8E",x"9C",x"5B",x"E6",x"86",x"0D",x"D8", -- 0x9B00
    x"27",x"18",x"BD",x"9B",x"98",x"81",x"23",x"27", -- 0x9B08
    x"04",x"81",x"2B",x"26",x"03",x"5C",x"20",x"0A", -- 0x9B10
    x"81",x"2D",x"26",x"03",x"5A",x"20",x"03",x"BD", -- 0x9B18
    x"9B",x"E2",x"5A",x"C1",x"0B",x"22",x"A6",x"34", -- 0x9B20
    x"04",x"D6",x"E1",x"96",x"E2",x"3D",x"DD",x"D5", -- 0x9B28
    x"33",x"61",x"96",x"DE",x"81",x"01",x"22",x"2C", -- 0x9B30
    x"8E",x"9C",x"62",x"C6",x"18",x"3D",x"3A",x"35", -- 0x9B38
    x"04",x"58",x"3A",x"31",x"84",x"8D",x"45",x"DD", -- 0x9B40
    x"E3",x"8D",x"0C",x"96",x"DF",x"8D",x"0B",x"8D", -- 0x9B48
    x"06",x"96",x"E0",x"8D",x"05",x"20",x"F2",x"86", -- 0x9B50
    x"7E",x"12",x"B7",x"FF",x"20",x"AE",x"A4",x"30", -- 0x9B58
    x"1F",x"26",x"FC",x"39",x"8E",x"9C",x"7A",x"C6", -- 0x9B60
    x"0C",x"3D",x"3A",x"35",x"04",x"3A",x"8D",x"1C", -- 0x9B68
    x"DD",x"E3",x"8D",x"0C",x"96",x"DF",x"8D",x"0B", -- 0x9B70
    x"8D",x"06",x"96",x"E0",x"8D",x"05",x"20",x"F2", -- 0x9B78
    x"86",x"7E",x"12",x"B7",x"FF",x"20",x"A6",x"84", -- 0x9B80
    x"4A",x"26",x"FD",x"39",x"C6",x"FF",x"96",x"E5", -- 0x9B88
    x"27",x"05",x"8B",x"02",x"3D",x"44",x"56",x"39", -- 0x9B90
    x"34",x"10",x"0D",x"D8",x"27",x"4D",x"9E",x"D9", -- 0x9B98
    x"A6",x"80",x"9F",x"D9",x"0A",x"D8",x"81",x"20", -- 0x9BA0
    x"27",x"F0",x"35",x"90",x"8D",x"EA",x"81",x"2B", -- 0x9BA8
    x"27",x"3C",x"81",x"2D",x"27",x"3C",x"81",x"3E", -- 0x9BB0
    x"27",x"42",x"81",x"3C",x"27",x"39",x"81",x"3D", -- 0x9BB8
    x"27",x"3F",x"BD",x"90",x"AA",x"25",x"24",x"5F", -- 0x9BC0
    x"80",x"30",x"97",x"D7",x"86",x"0A",x"3D",x"4D", -- 0x9BC8
    x"26",x"19",x"DB",x"D7",x"25",x"15",x"0D",x"D8", -- 0x9BD0
    x"27",x"17",x"BD",x"9B",x"98",x"BD",x"90",x"AA", -- 0x9BD8
    x"24",x"E6",x"0C",x"D8",x"9E",x"D9",x"30",x"1F", -- 0x9BE0
    x"9F",x"D9",x"39",x"7E",x"B4",x"4A",x"5C",x"27", -- 0x9BE8
    x"FA",x"39",x"5D",x"27",x"F6",x"5A",x"39",x"5D", -- 0x9BF0
    x"27",x"F1",x"54",x"39",x"5D",x"2B",x"EC",x"58", -- 0x9BF8
    x"39",x"34",x"60",x"8D",x"16",x"BD",x"B7",x"0E", -- 0x9C00
    x"35",x"E0",x"BD",x"9C",x"1B",x"C6",x"02",x"BD", -- 0x9C08
    x"AC",x"33",x"D6",x"D8",x"9E",x"D9",x"34",x"14", -- 0x9C10
    x"7E",x"9A",x"32",x"9E",x"D9",x"34",x"10",x"BD", -- 0x9C18
    x"9B",x"98",x"BD",x"B3",x"A2",x"25",x"C4",x"BD", -- 0x9C20
    x"9B",x"98",x"81",x"3B",x"26",x"F9",x"35",x"10", -- 0x9C28
    x"DE",x"A6",x"34",x"40",x"9F",x"A6",x"BD",x"B2", -- 0x9C30
    x"84",x"35",x"10",x"9F",x"A6",x"39",x"4F",x"1F", -- 0x9C38
    x"8B",x"DC",x"E3",x"10",x"27",x"0D",x"74",x"93", -- 0x9C40
    x"D5",x"DD",x"E3",x"22",x"0D",x"0F",x"E3",x"0F", -- 0x9C48
    x"E4",x"35",x"02",x"10",x"EE",x"67",x"84",x"7F", -- 0x9C50
    x"34",x"02",x"3B",x"0A",x"0C",x"01",x"03",x"05", -- 0x9C58
    x"06",x"08",x"01",x"A8",x"01",x"90",x"01",x"7A", -- 0x9C60
    x"01",x"64",x"01",x"50",x"01",x"3D",x"01",x"2B", -- 0x9C68
    x"01",x"1A",x"01",x"0A",x"00",x"FB",x"00",x"ED", -- 0x9C70
    x"00",x"DF",x"00",x"D3",x"00",x"C7",x"00",x"BB", -- 0x9C78
    x"00",x"B1",x"00",x"A6",x"00",x"9D",x"00",x"94", -- 0x9C80
    x"00",x"8B",x"00",x"83",x"00",x"7C",x"00",x"75", -- 0x9C88
    x"00",x"6E",x"A6",x"9C",x"93",x"8B",x"83",x"7B", -- 0x9C90
    x"74",x"6D",x"67",x"61",x"5B",x"56",x"51",x"4C", -- 0x9C98
    x"47",x"43",x"3F",x"3B",x"37",x"34",x"31",x"2E", -- 0x9CA0
    x"2B",x"28",x"26",x"23",x"21",x"1F",x"1D",x"1B", -- 0x9CA8
    x"19",x"18",x"16",x"14",x"13",x"12",x"9E",x"8A", -- 0x9CB0
    x"C6",x"01",x"34",x"14",x"D7",x"C2",x"9F",x"D5", -- 0x9CB8
    x"BD",x"95",x"9A",x"BD",x"B1",x"56",x"BD",x"B6", -- 0x9CC0
    x"54",x"20",x"08",x"BD",x"9B",x"98",x"7E",x"9B", -- 0x9CC8
    x"BE",x"35",x"14",x"D7",x"D8",x"27",x"FA",x"9F", -- 0x9CD0
    x"D9",x"10",x"27",x"00",x"EA",x"0D",x"D8",x"27", -- 0x9CD8
    x"F0",x"BD",x"9B",x"98",x"81",x"3B",x"27",x"F5", -- 0x9CE0
    x"81",x"27",x"27",x"F1",x"81",x"4E",x"26",x"04", -- 0x9CE8
    x"03",x"D5",x"20",x"E9",x"81",x"42",x"26",x"04", -- 0x9CF0
    x"03",x"D6",x"20",x"E1",x"81",x"58",x"10",x"27", -- 0x9CF8
    x"00",x"96",x"81",x"4D",x"10",x"27",x"01",x"2A", -- 0x9D00
    x"34",x"02",x"C6",x"01",x"0D",x"D8",x"27",x"11", -- 0x9D08
    x"BD",x"9B",x"98",x"BD",x"B3",x"A2",x"34",x"01", -- 0x9D10
    x"BD",x"9B",x"E2",x"35",x"01",x"24",x"02",x"8D", -- 0x9D18
    x"AA",x"35",x"02",x"81",x"43",x"27",x"28",x"81", -- 0x9D20
    x"41",x"27",x"2E",x"81",x"53",x"27",x"32",x"81", -- 0x9D28
    x"55",x"27",x"5C",x"81",x"44",x"27",x"55",x"81", -- 0x9D30
    x"4C",x"27",x"4C",x"81",x"52",x"27",x"43",x"80", -- 0x9D38
    x"45",x"27",x"2F",x"4A",x"27",x"27",x"4A",x"27", -- 0x9D40
    x"32",x"4A",x"27",x"1D",x"7E",x"B4",x"4A",x"BD", -- 0x9D48
    x"95",x"5D",x"D7",x"B2",x"BD",x"95",x"9A",x"20", -- 0x9D50
    x"84",x"C1",x"04",x"24",x"EF",x"D7",x"E8",x"20", -- 0x9D58
    x"F6",x"C1",x"3F",x"24",x"E7",x"D7",x"E9",x"20", -- 0x9D60
    x"EE",x"4F",x"8D",x"58",x"21",x"4F",x"1F",x"01", -- 0x9D68
    x"20",x"59",x"4F",x"1F",x"01",x"8D",x"4D",x"1E", -- 0x9D70
    x"01",x"20",x"50",x"4F",x"1F",x"01",x"8D",x"44", -- 0x9D78
    x"20",x"49",x"4F",x"9E",x"8A",x"20",x"44",x"4F", -- 0x9D80
    x"8D",x"3A",x"20",x"F7",x"4F",x"20",x"03",x"4F", -- 0x9D88
    x"8D",x"32",x"9E",x"8A",x"1E",x"10",x"20",x"33", -- 0x9D90
    x"BD",x"9C",x"1B",x"C6",x"02",x"BD",x"AC",x"33", -- 0x9D98
    x"D6",x"D8",x"9E",x"D9",x"34",x"14",x"7E",x"9C", -- 0x9DA0
    x"C6",x"D6",x"E9",x"27",x"1B",x"4F",x"1E",x"01", -- 0x9DA8
    x"A7",x"E2",x"2A",x"02",x"8D",x"0D",x"BD",x"9F", -- 0x9DB0
    x"B5",x"1F",x"30",x"44",x"56",x"44",x"56",x"6D", -- 0x9DB8
    x"E0",x"2A",x"04",x"40",x"50",x"82",x"00",x"39", -- 0x9DC0
    x"1F",x"10",x"39",x"34",x"06",x"8D",x"DA",x"35", -- 0x9DC8
    x"10",x"34",x"06",x"8D",x"D4",x"35",x"10",x"10", -- 0x9DD0
    x"9E",x"E8",x"34",x"20",x"6D",x"E4",x"27",x"08", -- 0x9DD8
    x"1E",x"10",x"8D",x"DF",x"6A",x"E4",x"20",x"F4", -- 0x9DE0
    x"35",x"20",x"DE",x"8A",x"D3",x"C7",x"2B",x"02", -- 0x9DE8
    x"1F",x"03",x"1F",x"10",x"9E",x"8A",x"D3",x"C9", -- 0x9DF0
    x"2B",x"02",x"1F",x"01",x"11",x"83",x"01",x"00", -- 0x9DF8
    x"25",x"03",x"CE",x"00",x"FF",x"8C",x"00",x"C0", -- 0x9E00
    x"25",x"03",x"8E",x"00",x"BF",x"DC",x"C7",x"DD", -- 0x9E08
    x"BD",x"DC",x"C9",x"DD",x"BF",x"9F",x"C5",x"DF", -- 0x9E10
    x"C3",x"0D",x"D5",x"26",x"04",x"9F",x"C9",x"DF", -- 0x9E18
    x"C7",x"BD",x"94",x"20",x"0D",x"D6",x"26",x"03", -- 0x9E20
    x"BD",x"94",x"A1",x"0F",x"D5",x"0F",x"D6",x"7E", -- 0x9E28
    x"9C",x"DD",x"BD",x"9B",x"98",x"34",x"02",x"BD", -- 0x9E30
    x"9E",x"5E",x"34",x"06",x"BD",x"9B",x"98",x"81", -- 0x9E38
    x"2C",x"10",x"26",x"FF",x"07",x"BD",x"9E",x"5B", -- 0x9E40
    x"1F",x"01",x"35",x"40",x"35",x"02",x"81",x"2B", -- 0x9E48
    x"27",x"04",x"81",x"2D",x"26",x"A6",x"1F",x"30", -- 0x9E50
    x"7E",x"9D",x"CB",x"BD",x"9B",x"98",x"81",x"2B", -- 0x9E58
    x"27",x"07",x"81",x"2D",x"27",x"04",x"BD",x"9B", -- 0x9E60
    x"E2",x"4F",x"34",x"02",x"BD",x"9C",x"CB",x"35", -- 0x9E68
    x"02",x"4D",x"27",x"04",x"4F",x"50",x"82",x"00", -- 0x9E70
    x"39",x"00",x"00",x"00",x"01",x"FE",x"C5",x"19", -- 0x9E78
    x"19",x"FB",x"16",x"31",x"F2",x"F4",x"FB",x"4A", -- 0x9E80
    x"51",x"EC",x"84",x"61",x"F9",x"E1",x"C7",x"78", -- 0x9E88
    x"AE",x"D4",x"DC",x"8E",x"3B",x"C5",x"E5",x"A2", -- 0x9E90
    x"69",x"B5",x"06",x"B5",x"06",x"81",x"40",x"26", -- 0x9E98
    x"02",x"9D",x"9F",x"BD",x"95",x"22",x"BD",x"93", -- 0x9EA0
    x"B2",x"BD",x"93",x"1D",x"AE",x"C4",x"9F",x"CB", -- 0x9EA8
    x"AE",x"42",x"9F",x"CD",x"BD",x"B2",x"6D",x"BD", -- 0x9EB0
    x"B7",x"3D",x"CE",x"00",x"CF",x"AF",x"C4",x"BD", -- 0x9EB8
    x"93",x"20",x"86",x"01",x"97",x"C2",x"BD",x"95", -- 0x9EC0
    x"81",x"8E",x"01",x"00",x"9D",x"A5",x"27",x"0F", -- 0x9EC8
    x"BD",x"B2",x"6D",x"BD",x"B1",x"41",x"96",x"4F", -- 0x9ED0
    x"8B",x"08",x"97",x"4F",x"BD",x"B7",x"40",x"96", -- 0x9ED8
    x"B6",x"85",x"02",x"27",x"04",x"1F",x"10",x"30", -- 0x9EE0
    x"8B",x"9F",x"D1",x"C6",x"01",x"D7",x"C2",x"D7", -- 0x9EE8
    x"D8",x"BD",x"9F",x"E2",x"34",x"06",x"BD",x"9F", -- 0x9EF0
    x"E2",x"DD",x"D9",x"35",x"06",x"34",x"06",x"9E", -- 0x9EF8
    x"11",x"3F",x"0F",x"03",x"CC",x"26",x"00",x"34", -- 0x9F00
    x"06",x"BE",x"C0",x"06",x"0C",x"03",x"96",x"03", -- 0x9F08
    x"81",x"12",x"22",x"22",x"A7",x"03",x"CC",x"02", -- 0x9F10
    x"00",x"A7",x"84",x"86",x"22",x"A7",x"02",x"35", -- 0x9F18
    x"06",x"ED",x"04",x"8B",x"01",x"34",x"06",x"AD", -- 0x9F20
    x"9F",x"C0",x"04",x"6D",x"06",x"27",x"DA",x"35", -- 0x9F28
    x"06",x"C6",x"28",x"7E",x"AC",x"46",x"35",x"06", -- 0x9F30
    x"FC",x"26",x"00",x"10",x"83",x"4F",x"53",x"10", -- 0x9F38
    x"27",x"46",x"BF",x"7F",x"26",x"00",x"7F",x"26", -- 0x9F40
    x"01",x"7E",x"A0",x"E8",x"CC",x"3B",x"3B",x"FD", -- 0x9F48
    x"01",x"00",x"FD",x"01",x"02",x"FD",x"01",x"04", -- 0x9F50
    x"39",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x9F58
    x"05",x"10",x"93",x"D3",x"25",x"02",x"DC",x"D3", -- 0x9F60
    x"DD",x"C3",x"A6",x"E4",x"81",x"04",x"25",x"0A", -- 0x9F68
    x"DC",x"CD",x"93",x"C5",x"24",x"11",x"4F",x"5F", -- 0x9F70
    x"20",x"0D",x"DC",x"CD",x"D3",x"C5",x"25",x"05", -- 0x9F78
    x"10",x"93",x"D5",x"25",x"02",x"DC",x"D5",x"DD", -- 0x9F80
    x"C5",x"0D",x"D8",x"26",x"02",x"8D",x"50",x"35", -- 0x9F88
    x"06",x"04",x"D8",x"25",x"05",x"10",x"93",x"D9", -- 0x9F90
    x"27",x"0C",x"5C",x"C1",x"08",x"26",x"04",x"4C", -- 0x9F98
    x"5F",x"84",x"07",x"7E",x"9E",x"FD",x"39",x"9E", -- 0x9FA0
    x"CF",x"EC",x"C4",x"27",x"07",x"83",x"00",x"01", -- 0x9FA8
    x"8D",x"03",x"1F",x"21",x"39",x"34",x"76",x"6F", -- 0x9FB0
    x"64",x"A6",x"63",x"3D",x"ED",x"66",x"EC",x"61", -- 0x9FB8
    x"3D",x"EB",x"66",x"89",x"00",x"ED",x"65",x"E6", -- 0x9FC0
    x"E4",x"A6",x"63",x"3D",x"E3",x"65",x"ED",x"65", -- 0x9FC8
    x"24",x"02",x"6C",x"64",x"A6",x"E4",x"E6",x"62", -- 0x9FD0
    x"3D",x"E3",x"64",x"ED",x"64",x"35",x"F6",x"7E", -- 0x9FD8
    x"94",x"A1",x"5F",x"9D",x"A5",x"27",x"11",x"BD", -- 0x9FE0
    x"B2",x"6D",x"BD",x"B1",x"41",x"96",x"4F",x"8B", -- 0x9FE8
    x"06",x"97",x"4F",x"BD",x"B7",x"0E",x"C4",x"3F", -- 0x9FF0
    x"1F",x"98",x"C4",x"07",x"44",x"44",x"44",x"39", -- 0x9FF8
    x"10",x"CE",x"00",x"FA",x"BD",x"DF",x"21",x"4F", -- 0xA000
    x"52",x"43",x"48",x"45",x"53",x"54",x"52",x"41", -- 0xA008
    x"2D",x"39",x"30",x"2F",x"43",x"43",x"20",x"28", -- 0xA010
    x"54",x"4D",x"29",x"0D",x"53",x"4F",x"46",x"54", -- 0xA018
    x"57",x"41",x"52",x"45",x"20",x"41",x"46",x"46", -- 0xA020
    x"41",x"49",x"52",x"2C",x"20",x"4C",x"54",x"44", -- 0xA028
    x"2E",x"0D",x"43",x"4F",x"50",x"59",x"52",x"49", -- 0xA030
    x"47",x"48",x"54",x"20",x"31",x"39",x"38",x"34", -- 0xA038
    x"20",x"4A",x"4F",x"4E",x"20",x"42",x"4F",x"4B", -- 0xA040
    x"45",x"4C",x"4D",x"41",x"4E",x"0D",x"4C",x"49", -- 0xA048
    x"43",x"45",x"4E",x"53",x"45",x"44",x"20",x"54", -- 0xA050
    x"4F",x"20",x"54",x"41",x"4E",x"44",x"59",x"20", -- 0xA058
    x"43",x"4F",x"52",x"50",x"4F",x"52",x"41",x"54", -- 0xA060
    x"49",x"4F",x"4E",x"0D",x"41",x"4C",x"4C",x"20", -- 0xA068
    x"52",x"49",x"47",x"48",x"54",x"53",x"20",x"52", -- 0xA070
    x"45",x"53",x"45",x"52",x"56",x"45",x"44",x"0D", -- 0xA078
    x"56",x"45",x"52",x"53",x"49",x"4F",x"4E",x"20", -- 0xA080
    x"30",x"31",x"2E",x"30",x"31",x"2E",x"30",x"30", -- 0xA088
    x"AF",x"20",x"57",x"49",x"4C",x"4C",x"49",x"41", -- 0xA090
    x"4D",x"20",x"54",x"45",x"4C",x"4C",x"20",x"4F", -- 0xA098
    x"56",x"45",x"52",x"54",x"55",x"52",x"45",x"AF", -- 0xA0A0
    x"20",x"42",x"59",x"20",x"52",x"4F",x"53",x"53", -- 0xA0A8
    x"49",x"4E",x"49",x"A0",x"A0",x"A0",x"A0",x"A0", -- 0xA0B0
    x"A0",x"CE",x"51",x"3D",x"36",x"36",x"5A",x"32", -- 0xA0B8
    x"4B",x"34",x"23",x"3C",x"33",x"4F",x"31",x"CD", -- 0xA0C0
    x"D9",x"41",x"28",x"51",x"2E",x"36",x"2C",x"53", -- 0xA0C8
    x"36",x"3B",x"36",x"3B",x"29",x"31",x"49",x"36", -- 0xA0D0
    x"3B",x"34",x"3B",x"32",x"3B",x"34",x"3B",x"36", -- 0xA0D8
    x"3B",x"34",x"3B",x"36",x"3B",x"39",x"3B",x"CD", -- 0xA0E0
    x"B6",x"3B",x"34",x"3B",x"32",x"3B",x"34",x"3B", -- 0xA0E8
    x"36",x"3B",x"34",x"3B",x"36",x"3B",x"39",x"3B", -- 0xA0F0
    x"D6",x"32",x"59",x"41",x"51",x"2E",x"32",x"2C", -- 0xA0F8
    x"53",x"32",x"3B",x"32",x"3B",x"51",x"2E",x"32", -- 0xA100
    x"2C",x"53",x"34",x"3B",x"34",x"3B",x"D6",x"33", -- 0xA108
    x"59",x"45",x"48",x"2E",x"2E",x"24",x"53",x"32", -- 0xA110
    x"3B",x"32",x"3B",x"CD",x"A8",x"51",x"2E",x"36", -- 0xA118
    x"2C",x"53",x"36",x"3B",x"36",x"3B",x"29",x"33", -- 0xA120
    x"D6",x"32",x"49",x"34",x"3B",x"33",x"3B",x"32", -- 0xA128
    x"3B",x"33",x"3B",x"34",x"3B",x"36",x"3B",x"35", -- 0xA130
    x"3B",x"34",x"3B",x"33",x"3B",x"34",x"3B",x"33", -- 0xA138
    x"3B",x"35",x"3B",x"34",x"3B",x"33",x"3B",x"32", -- 0xA140
    x"3B",x"34",x"3B",x"D6",x"33",x"32",x"3B",x"40", -- 0xA148
    x"31",x"3B",x"33",x"3B",x"31",x"3B",x"2A",x"32", -- 0xA150
    x"3B",x"34",x"3B",x"33",x"3B",x"32",x"3B",x"2D", -- 0xA158
    x"31",x"3B",x"32",x"3B",x"2D",x"31",x"3B",x"33", -- 0xA160
    x"3B",x"32",x"3B",x"2D",x"31",x"3B",x"2D",x"33", -- 0xA168
    x"3B",x"32",x"3B",x"D0",x"30",x"33",x"B6",x"3B", -- 0xA170
    x"53",x"28",x"36",x"3B",x"36",x"3B",x"49",x"29", -- 0xA178
    x"31",x"D6",x"32",x"33",x"3B",x"53",x"28",x"33", -- 0xA180
    x"3B",x"33",x"3B",x"49",x"29",x"31",x"D6",x"33", -- 0xA188
    x"28",x"31",x"3B",x"53",x"31",x"3B",x"31",x"3B", -- 0xA190
    x"49",x"31",x"3B",x"31",x"3B",x"C0",x"56",x"34", -- 0xA198
    x"59",x"41",x"29",x"31",x"A8",x"52",x"30",x"33", -- 0xA1A0
    x"29",x"32",x"D0",x"20",x"AA",x"57",x"36",x"D6", -- 0xA1A8
    x"32",x"33",x"D6",x"33",x"31",x"C0",x"56",x"34", -- 0xA1B0
    x"46",x"48",x"24",x"D0",x"30",x"35",x"D5",x"2B", -- 0xA1B8
    x"37",x"53",x"31",x"3B",x"31",x"3B",x"D6",x"33", -- 0xA1C0
    x"59",x"42",x"33",x"3B",x"33",x"3B",x"D6",x"34", -- 0xA1C8
    x"35",x"3B",x"35",x"3B",x"D0",x"30",x"36",x"A8", -- 0xA1D0
    x"4D",x"B1",x"31",x"2C",x"31",x"3B",x"31",x"3B", -- 0xA1D8
    x"D6",x"33",x"33",x"33",x"2C",x"33",x"3B",x"33", -- 0xA1E0
    x"3B",x"D6",x"34",x"35",x"35",x"2C",x"35",x"3B", -- 0xA1E8
    x"35",x"3B",x"29",x"31",x"D0",x"30",x"37",x"AA", -- 0xA1F0
    x"49",x"32",x"2C",x"33",x"2C",x"34",x"2C",x"40", -- 0xA1F8
    x"53",x"31",x"3B",x"31",x"3B",x"D6",x"32",x"49", -- 0xA200
    x"28",x"31",x"2C",x"29",x"32",x"D6",x"33",x"28", -- 0xA208
    x"33",x"2C",x"29",x"32",x"53",x"33",x"3B",x"33", -- 0xA210
    x"3B",x"D6",x"34",x"49",x"28",x"35",x"2C",x"29", -- 0xA218
    x"32",x"53",x"35",x"3B",x"35",x"3B",x"CD",x"B1", -- 0xA220
    x"31",x"2C",x"31",x"3B",x"31",x"3B",x"2A",x"32", -- 0xA228
    x"32",x"2C",x"34",x"3B",x"34",x"3B",x"C0",x"56", -- 0xA230
    x"32",x"51",x"24",x"49",x"28",x"31",x"3B",x"53", -- 0xA238
    x"29",x"32",x"A8",x"56",x"33",x"33",x"33",x"2C", -- 0xA240
    x"33",x"3B",x"33",x"3B",x"D6",x"34",x"35",x"35", -- 0xA248
    x"2C",x"35",x"3B",x"35",x"3B",x"29",x"31",x"CD", -- 0xA250
    x"AA",x"49",x"33",x"2C",x"31",x"2C",x"40",x"31", -- 0xA258
    x"2C",x"53",x"31",x"3B",x"31",x"3B",x"D6",x"32", -- 0xA260
    x"49",x"28",x"31",x"2C",x"29",x"32",x"D6",x"33", -- 0xA268
    x"28",x"34",x"2C",x"29",x"32",x"53",x"33",x"3B", -- 0xA270
    x"33",x"3B",x"D6",x"34",x"49",x"28",x"36",x"2C", -- 0xA278
    x"29",x"32",x"53",x"35",x"3B",x"35",x"3B",x"D2", -- 0xA280
    x"30",x"36",x"D0",x"30",x"38",x"AA",x"49",x"32", -- 0xA288
    x"2C",x"33",x"2C",x"34",x"2C",x"53",x"32",x"34", -- 0xA290
    x"C0",x"56",x"32",x"49",x"28",x"31",x"2C",x"29", -- 0xA298
    x"32",x"53",x"31",x"3B",x"31",x"3B",x"D6",x"33", -- 0xA2A0
    x"49",x"28",x"33",x"2C",x"29",x"32",x"53",x"33", -- 0xA2A8
    x"3B",x"33",x"3B",x"D6",x"34",x"49",x"28",x"35", -- 0xA2B0
    x"2C",x"29",x"32",x"53",x"35",x"3B",x"35",x"3B", -- 0xA2B8
    x"CD",x"AA",x"51",x"36",x"53",x"36",x"35",x"34", -- 0xA2C0
    x"33",x"C0",x"28",x"56",x"32",x"32",x"32",x"2C", -- 0xA2C8
    x"32",x"3B",x"32",x"3B",x"D6",x"33",x"36",x"36", -- 0xA2D0
    x"2C",x"36",x"3B",x"36",x"3B",x"D6",x"34",x"38", -- 0xA2D8
    x"38",x"2C",x"38",x"3B",x"38",x"3B",x"29",x"31", -- 0xA2E0
    x"CD",x"AA",x"49",x"32",x"3B",x"34",x"3B",x"32", -- 0xA2E8
    x"3B",x"C0",x"56",x"32",x"24",x"31",x"3B",x"31", -- 0xA2F0
    x"3B",x"A8",x"56",x"33",x"33",x"3B",x"D6",x"34", -- 0xA2F8
    x"35",x"3B",x"29",x"32",x"D2",x"30",x"35",x"59", -- 0xA300
    x"45",x"56",x"33",x"59",x"45",x"52",x"30",x"36", -- 0xA308
    x"52",x"30",x"37",x"52",x"30",x"36",x"52",x"30", -- 0xA310
    x"38",x"D0",x"20",x"AA",x"55",x"30",x"59",x"41", -- 0xA318
    x"53",x"42",x"3B",x"42",x"3B",x"D6",x"32",x"39", -- 0xA320
    x"3B",x"39",x"3B",x"C0",x"56",x"33",x"59",x"41", -- 0xA328
    x"30",x"3B",x"30",x"3B",x"D6",x"34",x"37",x"3B", -- 0xA330
    x"37",x"3B",x"D0",x"31",x"33",x"A8",x"4D",x"AA", -- 0xA338
    x"42",x"42",x"2C",x"42",x"3B",x"42",x"3B",x"D6", -- 0xA340
    x"32",x"39",x"39",x"2C",x"39",x"3B",x"39",x"3B", -- 0xA348
    x"D6",x"33",x"30",x"30",x"2C",x"30",x"3B",x"30", -- 0xA350
    x"3B",x"C0",x"56",x"34",x"37",x"37",x"2C",x"37", -- 0xA358
    x"3B",x"37",x"3B",x"29",x"31",x"A8",x"4D",x"AA", -- 0xA360
    x"49",x"42",x"3B",x"45",x"3B",x"D6",x"32",x"39", -- 0xA368
    x"3B",x"37",x"3B",x"D6",x"33",x"30",x"3B",x"24", -- 0xA370
    x"D6",x"34",x"2D",x"37",x"3B",x"24",x"29",x"31", -- 0xA378
    x"D0",x"31",x"34",x"C2",x"3B",x"45",x"3B",x"42", -- 0xA380
    x"3B",x"41",x"3B",x"39",x"3B",x"38",x"3B",x"37", -- 0xA388
    x"3B",x"53",x"42",x"3B",x"42",x"3B",x"D6",x"32", -- 0xA390
    x"49",x"39",x"3B",x"37",x"3B",x"39",x"3B",x"38", -- 0xA398
    x"3B",x"37",x"3B",x"37",x"3B",x"34",x"3B",x"53", -- 0xA3A0
    x"39",x"3B",x"39",x"3B",x"C0",x"56",x"33",x"49", -- 0xA3A8
    x"30",x"3B",x"24",x"33",x"3B",x"24",x"33",x"3B", -- 0xA3B0
    x"34",x"3B",x"35",x"3B",x"53",x"30",x"3B",x"30", -- 0xA3B8
    x"3B",x"D6",x"34",x"49",x"37",x"3B",x"24",x"41", -- 0xA3C0
    x"3B",x"24",x"28",x"37",x"3B",x"29",x"32",x"53", -- 0xA3C8
    x"37",x"3B",x"37",x"3B",x"D2",x"31",x"33",x"D0", -- 0xA3D0
    x"31",x"35",x"AA",x"49",x"42",x"3B",x"45",x"3B", -- 0xA3D8
    x"44",x"3B",x"43",x"23",x"3B",x"D6",x"32",x"39", -- 0xA3E0
    x"3B",x"37",x"3B",x"41",x"3B",x"39",x"3B",x"D6", -- 0xA3E8
    x"33",x"30",x"3B",x"24",x"31",x"3B",x"30",x"3B", -- 0xA3F0
    x"C0",x"56",x"34",x"37",x"3B",x"24",x"34",x"3B", -- 0xA3F8
    x"34",x"3B",x"D0",x"20",x"AA",x"44",x"3B",x"43", -- 0xA400
    x"23",x"3B",x"44",x"3B",x"53",x"42",x"23",x"3B", -- 0xA408
    x"42",x"3B",x"D6",x"32",x"49",x"38",x"3B",x"37", -- 0xA410
    x"3B",x"38",x"3B",x"53",x"39",x"3B",x"39",x"3B", -- 0xA418
    x"C0",x"56",x"33",x"49",x"31",x"3B",x"32",x"23", -- 0xA420
    x"3B",x"31",x"3B",x"53",x"30",x"3B",x"30",x"3B", -- 0xA428
    x"D6",x"34",x"49",x"28",x"38",x"3B",x"29",x"32", -- 0xA430
    x"53",x"37",x"3B",x"37",x"3B",x"D2",x"31",x"33", -- 0xA438
    x"52",x"31",x"34",x"52",x"31",x"33",x"52",x"31", -- 0xA440
    x"35",x"D0",x"20",x"AA",x"28",x"44",x"3B",x"43", -- 0xA448
    x"23",x"3B",x"45",x"3B",x"43",x"3B",x"29",x"33", -- 0xA450
    x"D6",x"32",x"38",x"3B",x"D6",x"33",x"59",x"43", -- 0xA458
    x"49",x"2D",x"31",x"3B",x"24",x"24",x"28",x"53", -- 0xA460
    x"33",x"3B",x"33",x"3B",x"49",x"33",x"3B",x"29", -- 0xA468
    x"31",x"34",x"3B",x"C0",x"56",x"34",x"38",x"3B", -- 0xA470
    x"24",x"24",x"28",x"53",x"31",x"3B",x"31",x"3B", -- 0xA478
    x"31",x"31",x"2C",x"29",x"31",x"2A",x"32",x"3B", -- 0xA480
    x"CD",x"A8",x"44",x"3B",x"43",x"23",x"3B",x"45", -- 0xA488
    x"3B",x"43",x"3B",x"29",x"33",x"D6",x"33",x"49", -- 0xA490
    x"35",x"3B",x"33",x"33",x"22",x"35",x"3B",x"34", -- 0xA498
    x"3B",x"32",x"32",x"22",x"34",x"3B",x"D6",x"34", -- 0xA4A0
    x"33",x"3B",x"2D",x"31",x"2D",x"31",x"22",x"33", -- 0xA4A8
    x"3B",x"32",x"3B",x"2D",x"33",x"2D",x"33",x"22", -- 0xA4B0
    x"32",x"3B",x"CD",x"D3",x"44",x"3B",x"43",x"23", -- 0xA4B8
    x"3B",x"45",x"3B",x"43",x"3B",x"49",x"44",x"2C", -- 0xA4C0
    x"C0",x"56",x"32",x"24",x"31",x"3B",x"31",x"3B", -- 0xA4C8
    x"D6",x"33",x"24",x"34",x"3B",x"34",x"3B",x"D6", -- 0xA4D0
    x"34",x"2B",x"33",x"3B",x"36",x"3B",x"36",x"3B", -- 0xA4D8
    x"D0",x"20",x"A8",x"4D",x"AA",x"59",x"42",x"53", -- 0xA4E0
    x"41",x"3B",x"41",x"3B",x"41",x"41",x"2C",x"D6", -- 0xA4E8
    x"32",x"59",x"43",x"36",x"3B",x"36",x"3B",x"36", -- 0xA4F0
    x"36",x"2C",x"D6",x"33",x"33",x"3B",x"33",x"3B", -- 0xA4F8
    x"33",x"33",x"2C",x"C0",x"56",x"34",x"31",x"3B", -- 0xA500
    x"31",x"3B",x"49",x"31",x"3B",x"29",x"31",x"CD", -- 0xA508
    x"AA",x"42",x"3B",x"43",x"2C",x"41",x"41",x"22", -- 0xA510
    x"43",x"3B",x"42",x"2C",x"39",x"39",x"22",x"42", -- 0xA518
    x"3B",x"41",x"2C",x"53",x"36",x"3B",x"36",x"3B", -- 0xA520
    x"49",x"36",x"3B",x"D6",x"32",x"39",x"3B",x"41", -- 0xA528
    x"2C",x"36",x"36",x"22",x"41",x"3B",x"39",x"2C", -- 0xA530
    x"34",x"34",x"22",x"39",x"3B",x"38",x"2C",x"D6", -- 0xA538
    x"34",x"32",x"3B",x"D6",x"33",x"34",x"3B",x"40", -- 0xA540
    x"28",x"2B",x"35",x"2C",x"38",x"2C",x"37",x"2C", -- 0xA548
    x"36",x"2C",x"35",x"2C",x"34",x"2C",x"33",x"2C", -- 0xA550
    x"32",x"2C",x"31",x"2C",x"D6",x"34",x"29",x"31", -- 0xA558
    x"D2",x"30",x"35",x"59",x"41",x"56",x"32",x"59", -- 0xA560
    x"41",x"56",x"33",x"59",x"41",x"52",x"30",x"36", -- 0xA568
    x"52",x"30",x"37",x"52",x"30",x"36",x"52",x"30", -- 0xA570
    x"38",x"D2",x"30",x"35",x"59",x"45",x"56",x"33", -- 0xA578
    x"59",x"45",x"52",x"30",x"36",x"52",x"30",x"37", -- 0xA580
    x"52",x"30",x"36",x"52",x"30",x"38",x"D0",x"20", -- 0xA588
    x"5A",x"31",x"AA",x"59",x"41",x"53",x"28",x"36", -- 0xA590
    x"3B",x"36",x"3B",x"D6",x"32",x"29",x"31",x"C0", -- 0xA598
    x"56",x"34",x"31",x"3B",x"31",x"3B",x"A8",x"4D", -- 0xA5A0
    x"AA",x"36",x"36",x"2C",x"36",x"3B",x"36",x"3B", -- 0xA5A8
    x"D6",x"32",x"36",x"36",x"2C",x"36",x"3B",x"36", -- 0xA5B0
    x"3B",x"C0",x"56",x"34",x"31",x"31",x"2C",x"31", -- 0xA5B8
    x"3B",x"31",x"3B",x"29",x"31",x"CD",x"AA",x"49", -- 0xA5C0
    x"28",x"42",x"3B",x"43",x"3B",x"44",x"3B",x"24", -- 0xA5C8
    x"39",x"3B",x"41",x"3B",x"42",x"3B",x"D6",x"32", -- 0xA5D0
    x"29",x"31",x"D6",x"34",x"34",x"3B",x"35",x"3B", -- 0xA5D8
    x"36",x"3B",x"24",x"32",x"3B",x"33",x"3B",x"34", -- 0xA5E0
    x"3B",x"24",x"CD",x"C2",x"3B",x"43",x"3B",x"44", -- 0xA5E8
    x"3B",x"D6",x"32",x"34",x"3B",x"35",x"3B",x"36", -- 0xA5F0
    x"3B",x"C0",x"56",x"34",x"33",x"3B",x"32",x"3B", -- 0xA5F8
    x"31",x"3B",x"48",x"24",x"CD",x"AA",x"53",x"36", -- 0xA600
    x"36",x"23",x"37",x"38",x"25",x"38",x"23",x"39", -- 0xA608
    x"39",x"23",x"41",x"C0",x"28",x"56",x"32",x"53", -- 0xA610
    x"34",x"3B",x"31",x"3B",x"D6",x"33",x"59",x"41", -- 0xA618
    x"36",x"3B",x"24",x"D6",x"34",x"38",x"3B",x"24", -- 0xA620
    x"29",x"33",x"CD",x"AA",x"55",x"2B",x"37",x"53", -- 0xA628
    x"34",x"25",x"34",x"23",x"35",x"35",x"23",x"36", -- 0xA630
    x"36",x"23",x"37",x"38",x"C0",x"28",x"56",x"32", -- 0xA638
    x"53",x"34",x"3B",x"31",x"3B",x"D6",x"33",x"36", -- 0xA640
    x"3B",x"24",x"D6",x"34",x"38",x"3B",x"24",x"29", -- 0xA648
    x"33",x"A8",x"4D",x"AA",x"59",x"43",x"53",x"39", -- 0xA650
    x"38",x"41",x"38",x"D6",x"32",x"59",x"44",x"39", -- 0xA658
    x"38",x"41",x"38",x"C0",x"56",x"33",x"49",x"33", -- 0xA660
    x"3B",x"32",x"3B",x"D6",x"34",x"35",x"3B",x"38", -- 0xA668
    x"3B",x"29",x"37",x"CD",x"AA",x"55",x"30",x"47", -- 0xA670
    x"3B",x"53",x"28",x"47",x"39",x"29",x"32",x"C0", -- 0xA678
    x"56",x"32",x"59",x"41",x"51",x"24",x"53",x"28", -- 0xA680
    x"31",x"3B",x"2B",x"32",x"3B",x"29",x"31",x"D6", -- 0xA688
    x"33",x"59",x"45",x"49",x"33",x"3B",x"24",x"53", -- 0xA690
    x"33",x"3B",x"24",x"33",x"3B",x"D6",x"34",x"49", -- 0xA698
    x"35",x"3B",x"24",x"53",x"35",x"3B",x"24",x"35", -- 0xA6A0
    x"CD",x"AA",x"49",x"47",x"3B",x"53",x"28",x"44", -- 0xA6A8
    x"36",x"29",x"32",x"49",x"44",x"3B",x"53",x"28", -- 0xA6B0
    x"42",x"34",x"29",x"32",x"49",x"42",x"3B",x"53", -- 0xA6B8
    x"28",x"39",x"32",x"29",x"32",x"C0",x"56",x"32", -- 0xA6C0
    x"28",x"49",x"31",x"3B",x"53",x"31",x"3B",x"31", -- 0xA6C8
    x"3B",x"49",x"31",x"3B",x"2B",x"32",x"3B",x"29", -- 0xA6D0
    x"31",x"A8",x"56",x"33",x"33",x"3B",x"53",x"33", -- 0xA6D8
    x"3B",x"33",x"3B",x"49",x"33",x"3B",x"31",x"3B", -- 0xA6E0
    x"D6",x"34",x"35",x"3B",x"53",x"35",x"3B",x"35", -- 0xA6E8
    x"3B",x"49",x"35",x"3B",x"33",x"3B",x"29",x"32", -- 0xA6F0
    x"CD",x"AA",x"28",x"39",x"3B",x"53",x"39",x"3B", -- 0xA6F8
    x"39",x"3B",x"49",x"39",x"3B",x"39",x"3B",x"39", -- 0xA700
    x"3B",x"53",x"36",x"3B",x"36",x"3B",x"49",x"36", -- 0xA708
    x"3B",x"36",x"3B",x"36",x"3B",x"D6",x"32",x"29", -- 0xA710
    x"31",x"C0",x"56",x"33",x"33",x"3B",x"28",x"2B", -- 0xA718
    x"32",x"3B",x"29",x"33",x"28",x"31",x"3B",x"29", -- 0xA720
    x"33",x"D6",x"34",x"28",x"35",x"3B",x"29",x"34", -- 0xA728
    x"28",x"38",x"3B",x"29",x"33",x"CD",x"AA",x"28", -- 0xA730
    x"53",x"34",x"3B",x"34",x"3B",x"49",x"34",x"3B", -- 0xA738
    x"34",x"3B",x"34",x"3B",x"53",x"32",x"3B",x"32", -- 0xA740
    x"3B",x"49",x"32",x"3B",x"32",x"3B",x"D6",x"32", -- 0xA748
    x"29",x"31",x"C0",x"56",x"33",x"28",x"33",x"3B", -- 0xA750
    x"29",x"33",x"28",x"35",x"3B",x"29",x"32",x"D6", -- 0xA758
    x"34",x"28",x"41",x"3B",x"29",x"33",x"28",x"43", -- 0xA760
    x"3B",x"29",x"32",x"CD",x"A8",x"2A",x"56",x"31", -- 0xA768
    x"32",x"3B",x"2D",x"31",x"3B",x"D6",x"32",x"32", -- 0xA770
    x"3B",x"2D",x"31",x"3B",x"C0",x"56",x"33",x"35", -- 0xA778
    x"3B",x"38",x"3B",x"29",x"31",x"D6",x"34",x"55", -- 0xA780
    x"37",x"43",x"3B",x"38",x"3B",x"35",x"3B",x"38", -- 0xA788
    x"3B",x"CD",x"AA",x"28",x"34",x"3B",x"32",x"3B", -- 0xA790
    x"36",x"3B",x"34",x"3B",x"39",x"3B",x"36",x"3B", -- 0xA798
    x"42",x"3B",x"39",x"3B",x"44",x"3B",x"42",x"3B", -- 0xA7A0
    x"D6",x"32",x"29",x"31",x"C0",x"56",x"33",x"28", -- 0xA7A8
    x"33",x"3B",x"35",x"3B",x"31",x"3B",x"33",x"3B", -- 0xA7B0
    x"35",x"3B",x"38",x"3B",x"33",x"3B",x"35",x"3B", -- 0xA7B8
    x"31",x"3B",x"33",x"3B",x"D6",x"34",x"29",x"31", -- 0xA7C0
    x"CD",x"AA",x"51",x"2E",x"47",x"2C",x"53",x"47", -- 0xA7C8
    x"3B",x"47",x"3B",x"D6",x"32",x"51",x"2E",x"42", -- 0xA7D0
    x"2C",x"53",x"42",x"3B",x"42",x"3B",x"D6",x"33", -- 0xA7D8
    x"55",x"37",x"51",x"2E",x"39",x"2C",x"53",x"39", -- 0xA7E0
    x"3B",x"39",x"3B",x"D6",x"34",x"51",x"2E",x"32", -- 0xA7E8
    x"2C",x"53",x"32",x"3B",x"32",x"3B",x"CD",x"A8", -- 0xA7F0
    x"56",x"31",x"49",x"47",x"3B",x"D6",x"32",x"42", -- 0xA7F8
    x"3B",x"D6",x"33",x"39",x"3B",x"29",x"33",x"D6", -- 0xA800
    x"34",x"32",x"40",x"31",x"33",x"31",x"CD",x"AA", -- 0xA808
    x"51",x"2E",x"47",x"2C",x"53",x"24",x"47",x"3B", -- 0xA810
    x"51",x"2E",x"47",x"2C",x"53",x"24",x"39",x"3B", -- 0xA818
    x"57",x"39",x"D6",x"32",x"51",x"2E",x"42",x"2C", -- 0xA820
    x"53",x"24",x"42",x"3B",x"51",x"2E",x"42",x"2C", -- 0xA828
    x"53",x"24",x"2D",x"33",x"3B",x"57",x"2D",x"33", -- 0xA830
    x"D6",x"33",x"51",x"2E",x"39",x"2C",x"53",x"24", -- 0xA838
    x"36",x"3B",x"51",x"2E",x"36",x"2C",x"40",x"53", -- 0xA840
    x"24",x"31",x"3B",x"57",x"31",x"D6",x"34",x"51", -- 0xA848
    x"2E",x"35",x"2C",x"53",x"24",x"35",x"3B",x"51", -- 0xA850
    x"2E",x"35",x"2C",x"53",x"24",x"43",x"3B",x"57", -- 0xA858
    x"43",x"39",x"BD",x"D7",x"0D",x"2B",x"15",x"8E", -- 0xA860
    x"CF",x"E2",x"BD",x"D6",x"50",x"25",x"3E",x"97", -- 0xA868
    x"96",x"A6",x"41",x"80",x"57",x"27",x"02",x"86", -- 0xA870
    x"FF",x"43",x"97",x"97",x"86",x"FE",x"97",x"6F", -- 0xA878
    x"9E",x"60",x"6D",x"84",x"2A",x"04",x"86",x"0D", -- 0xA880
    x"8D",x"10",x"A6",x"80",x"84",x"7F",x"27",x"D1", -- 0xA888
    x"81",x"60",x"25",x"02",x"80",x"40",x"8D",x"02", -- 0xA890
    x"20",x"E8",x"6E",x"9F",x"A0",x"02",x"BD",x"CA", -- 0xA898
    x"DF",x"9E",x"62",x"69",x"84",x"4F",x"66",x"84", -- 0xA8A0
    x"BD",x"CA",x"C2",x"20",x"36",x"7E",x"CC",x"02", -- 0xA8A8
    x"C6",x"02",x"5A",x"D7",x"58",x"9E",x"62",x"96", -- 0xA8B0
    x"58",x"30",x"86",x"9C",x"74",x"22",x"EE",x"9C", -- 0xA8B8
    x"5E",x"25",x"EA",x"34",x"10",x"33",x"21",x"A6", -- 0xA8C0
    x"C0",x"2B",x"16",x"A8",x"80",x"48",x"27",x"F7", -- 0xA8C8
    x"35",x"10",x"20",x"E3",x"0D",x"B9",x"26",x"02", -- 0xA8D0
    x"0C",x"5C",x"10",x"AF",x"E4",x"8D",x"29",x"35", -- 0xA8D8
    x"90",x"35",x"10",x"9F",x"62",x"30",x"01",x"6D", -- 0xA8E0
    x"82",x"2A",x"FC",x"BD",x"CA",x"BB",x"33",x"88", -- 0xA8E8
    x"1E",x"11",x"93",x"62",x"24",x"40",x"A6",x"84", -- 0xA8F0
    x"48",x"27",x"39",x"C6",x"1F",x"30",x"01",x"6D", -- 0xA8F8
    x"84",x"2B",x"E8",x"5A",x"26",x"F7",x"20",x"E3", -- 0xA900
    x"8E",x"04",x"20",x"20",x"0C",x"9E",x"74",x"9F", -- 0xA908
    x"5D",x"9F",x"5E",x"7E",x"CA",x"B9",x"8E",x"04", -- 0xA910
    x"00",x"86",x"01",x"C6",x"8F",x"E7",x"80",x"1E", -- 0xA918
    x"10",x"C5",x"1F",x"1E",x"10",x"26",x"F6",x"4A", -- 0xA920
    x"26",x"F3",x"39",x"9E",x"74",x"8D",x"E0",x"9E", -- 0xA928
    x"5E",x"8C",x"9E",x"74",x"8D",x"DD",x"86",x"06", -- 0xA930
    x"DE",x"60",x"C6",x"1F",x"11",x"93",x"5E",x"27", -- 0xA938
    x"0A",x"6D",x"C2",x"2B",x"03",x"5A",x"26",x"F9", -- 0xA940
    x"4A",x"26",x"EF",x"8E",x"04",x"40",x"E6",x"1F", -- 0xA948
    x"D7",x"6B",x"4D",x"27",x"02",x"8D",x"C4",x"30", -- 0xA950
    x"1F",x"D6",x"6B",x"F7",x"04",x"3F",x"1F",x"10", -- 0xA958
    x"CA",x"E0",x"5C",x"27",x"04",x"6D",x"C4",x"2A", -- 0xA960
    x"0B",x"69",x"C4",x"53",x"66",x"C4",x"8D",x"A9", -- 0xA968
    x"9C",x"AD",x"27",x"26",x"E6",x"C4",x"C4",x"7F", -- 0xA970
    x"26",x"02",x"C6",x"8F",x"11",x"93",x"62",x"26", -- 0xA978
    x"0C",x"9F",x"88",x"0D",x"55",x"26",x"06",x"C8", -- 0xA980
    x"40",x"2A",x"02",x"C8",x"4F",x"E7",x"80",x"E6", -- 0xA988
    x"C0",x"58",x"26",x"C5",x"8D",x"83",x"9C",x"AD", -- 0xA990
    x"26",x"FA",x"39",x"03",x"CB",x"E1",x"0A",x"CA", -- 0xA998
    x"84",x"0B",x"CA",x"70",x"0D",x"CA",x"80",x"1A", -- 0xA9A0
    x"CA",x"A7",x"1B",x"C8",x"9E",x"1D",x"CA",x"80", -- 0xA9A8
    x"21",x"CA",x"D1",x"3F",x"CA",x"7C",x"FF",x"A6", -- 0xA9B0
    x"01",x"A7",x"80",x"6D",x"84",x"2A",x"F8",x"39", -- 0xA9B8
    x"30",x"A8",x"1F",x"9C",x"88",x"27",x"06",x"A6", -- 0xA9C0
    x"82",x"A7",x"01",x"20",x"F6",x"86",x"60",x"A7", -- 0xA9C8
    x"84",x"39",x"03",x"DD",x"A4",x"08",x"CA",x"62", -- 0xA9D0
    x"09",x"CA",x"5B",x"0C",x"CB",x"2C",x"0D",x"C8", -- 0xA9D8
    x"DA",x"13",x"CA",x"12",x"18",x"C9",x"BB",x"19", -- 0xA9E0
    x"C9",x"C0",x"1C",x"CB",x"3C",x"1D",x"C8",x"D4", -- 0xA9E8
    x"FF",x"8E",x"00",x"53",x"C6",x"0A",x"6F",x"80", -- 0xA9F0
    x"5A",x"26",x"FB",x"39",x"10",x"8E",x"04",x"00", -- 0xA9F8
    x"0D",x"58",x"26",x"03",x"BD",x"C9",x"16",x"10", -- 0xAA00
    x"9F",x"88",x"8D",x"E5",x"20",x"14",x"BD",x"C9", -- 0xAA08
    x"16",x"5A",x"5C",x"D7",x"58",x"BD",x"C9",x"08", -- 0xAA10
    x"10",x"8E",x"05",x"00",x"C6",x"08",x"D7",x"55", -- 0xAA18
    x"D7",x"54",x"F7",x"FF",x"22",x"0D",x"54",x"27", -- 0xAA20
    x"03",x"BD",x"C9",x"36",x"C6",x"8F",x"E7",x"A8", -- 0xAA28
    x"1F",x"BD",x"CC",x"09",x"8D",x"02",x"20",x"ED", -- 0xAA30
    x"97",x"54",x"0D",x"55",x"27",x"06",x"8E",x"C9", -- 0xAA38
    x"9B",x"BD",x"CB",x"D1",x"0F",x"54",x"8E",x"C9", -- 0xAA40
    x"D2",x"BD",x"CB",x"D1",x"81",x"20",x"25",x"0A", -- 0xAA48
    x"8A",x"40",x"A7",x"80",x"1F",x"10",x"C5",x"20", -- 0xAA50
    x"27",x"13",x"39",x"6D",x"80",x"2A",x"0E",x"0F", -- 0xAA58
    x"89",x"39",x"0A",x"89",x"2A",x"FB",x"8C",x"30", -- 0xAA60
    x"01",x"6D",x"84",x"2A",x"FA",x"9F",x"88",x"39", -- 0xAA68
    x"8D",x"6D",x"9C",x"5E",x"27",x"1E",x"6D",x"82", -- 0xAA70
    x"2A",x"F8",x"20",x"18",x"9E",x"74",x"8D",x"39", -- 0xAA78
    x"1F",x"21",x"9F",x"88",x"8D",x"59",x"9C",x"74", -- 0xAA80
    x"27",x"2F",x"30",x"01",x"6D",x"84",x"2A",x"F6", -- 0xAA88
    x"9C",x"74",x"27",x"25",x"8D",x"25",x"5F",x"D1", -- 0xAA90
    x"89",x"27",x"06",x"5C",x"6D",x"85",x"2A",x"F7", -- 0xAA98
    x"5A",x"3A",x"9F",x"62",x"9E",x"60",x"39",x"8D", -- 0xAAA0
    x"36",x"9E",x"62",x"D6",x"89",x"26",x"0C",x"C6", -- 0xAAA8
    x"01",x"8D",x"5D",x"9E",x"62",x"C6",x"60",x"E7", -- 0xAAB0
    x"82",x"9F",x"62",x"9F",x"60",x"69",x"84",x"53", -- 0xAAB8
    x"66",x"84",x"C6",x"80",x"E7",x"9F",x"00",x"74", -- 0xAAC0
    x"EA",x"9F",x"00",x"5E",x"E7",x"9F",x"00",x"5E", -- 0xAAC8
    x"39",x"0F",x"89",x"8E",x"08",x"00",x"BD",x"C9", -- 0xAAD0
    x"19",x"8D",x"95",x"8D",x"CC",x"1F",x"21",x"1F", -- 0xAAD8
    x"10",x"5F",x"1F",x"01",x"5A",x"5C",x"6D",x"85", -- 0xAAE0
    x"2A",x"FB",x"34",x"06",x"4F",x"9E",x"60",x"9C", -- 0xAAE8
    x"74",x"27",x"07",x"4C",x"6D",x"86",x"2A",x"FB", -- 0xAAF0
    x"30",x"86",x"34",x"16",x"E0",x"E0",x"27",x"02", -- 0xAAF8
    x"8D",x"0E",x"35",x"54",x"5D",x"27",x"8D",x"A6", -- 0xAB00
    x"C2",x"A7",x"82",x"5A",x"26",x"F9",x"20",x"84", -- 0xAB08
    x"D7",x"5D",x"50",x"2A",x"36",x"9E",x"5E",x"33", -- 0xAB10
    x"85",x"11",x"83",x"10",x"64",x"10",x"23",x"06", -- 0xAB18
    x"F8",x"DF",x"5E",x"A6",x"80",x"A7",x"C0",x"9C", -- 0xAB20
    x"60",x"25",x"F8",x"39",x"BD",x"C9",x"19",x"0D", -- 0xAB28
    x"55",x"27",x"08",x"0D",x"89",x"26",x"04",x"C6", -- 0xAB30
    x"60",x"E7",x"A4",x"39",x"1F",x"21",x"9F",x"88", -- 0xAB38
    x"BD",x"C9",x"19",x"0D",x"55",x"27",x"F4",x"0C", -- 0xAB40
    x"54",x"20",x"94",x"9E",x"60",x"33",x"85",x"A6", -- 0xAB48
    x"82",x"A7",x"C2",x"9C",x"5E",x"22",x"F8",x"27", -- 0xAB50
    x"02",x"33",x"41",x"DF",x"5E",x"39",x"40",x"D4", -- 0xAB58
    x"8D",x"41",x"D1",x"70",x"42",x"C9",x"32",x"43", -- 0xAB60
    x"D0",x"21",x"44",x"D3",x"2D",x"45",x"CA",x"0E", -- 0xAB68
    x"47",x"CB",x"B9",x"4B",x"D2",x"F8",x"4C",x"C8", -- 0xAB70
    x"62",x"4D",x"CB",x"AA",x"4E",x"C9",x"2B",x"4F", -- 0xAB78
    x"DC",x"AC",x"50",x"D8",x"5B",x"52",x"D1",x"69", -- 0xAB80
    x"53",x"D4",x"B9",x"54",x"C9",x"2F",x"56",x"D1", -- 0xAB88
    x"62",x"57",x"D0",x"A8",x"58",x"DD",x"AB",x"61", -- 0xAB90
    x"DA",x"1F",x"6D",x"C8",x"B2",x"6F",x"C8",x"B0", -- 0xAB98
    x"74",x"D4",x"D3",x"75",x"D4",x"D3",x"7F",x"DA", -- 0xABA0
    x"23",x"FF",x"BD",x"D7",x"0D",x"2B",x"31",x"97", -- 0xABA8
    x"58",x"96",x"58",x"27",x"34",x"10",x"8E",x"04", -- 0xABB0
    x"00",x"10",x"9F",x"64",x"97",x"57",x"32",x"62", -- 0xABB8
    x"10",x"9E",x"64",x"BD",x"D1",x"69",x"BD",x"CE", -- 0xABC0
    x"B7",x"BD",x"D4",x"B9",x"BD",x"D8",x"69",x"20", -- 0xABC8
    x"EF",x"30",x"03",x"A1",x"1D",x"25",x"06",x"26", -- 0xABD0
    x"F8",x"AE",x"1E",x"AF",x"E4",x"9E",x"88",x"5F", -- 0xABD8
    x"39",x"BD",x"CA",x"DF",x"0F",x"55",x"BD",x"C9", -- 0xABE0
    x"36",x"10",x"CE",x"00",x"FA",x"BD",x"CE",x"B7", -- 0xABE8
    x"8D",x"02",x"20",x"F5",x"8D",x"65",x"BD",x"C9", -- 0xABF0
    x"FC",x"A6",x"A4",x"2B",x"EC",x"8E",x"CB",x"5E", -- 0xABF8
    x"8D",x"CF",x"CC",x"7F",x"7F",x"FD",x"04",x"20", -- 0xAC00
    x"39",x"0F",x"6A",x"9E",x"88",x"E6",x"84",x"D7", -- 0xAC08
    x"AF",x"8D",x"0C",x"0D",x"B0",x"27",x"FA",x"96", -- 0xAC10
    x"87",x"08",x"94",x"25",x"F4",x"20",x"25",x"9E", -- 0xAC18
    x"88",x"E6",x"84",x"0D",x"6A",x"26",x"06",x"C8", -- 0xAC20
    x"40",x"2A",x"02",x"C8",x"4F",x"E7",x"84",x"8D", -- 0xAC28
    x"2A",x"26",x"09",x"0A",x"6A",x"D6",x"6A",x"C5", -- 0xAC30
    x"3F",x"26",x"E4",x"39",x"32",x"62",x"97",x"87", -- 0xAC38
    x"C6",x"FC",x"D7",x"94",x"D6",x"AF",x"E7",x"9F", -- 0xAC40
    x"00",x"88",x"39",x"8E",x"04",x"5E",x"0D",x"70", -- 0xAC48
    x"10",x"27",x"07",x"B4",x"C6",x"9D",x"13",x"5A", -- 0xAC50
    x"26",x"FC",x"39",x"CE",x"FF",x"00",x"8E",x"00", -- 0xAC58
    x"B0",x"6F",x"80",x"4F",x"4A",x"34",x"12",x"A7", -- 0xAC60
    x"42",x"69",x"42",x"24",x"3E",x"6C",x"E4",x"8D", -- 0xAC68
    x"7B",x"A7",x"61",x"1F",x"89",x"A8",x"84",x"E7", -- 0xAC70
    x"84",x"DA",x"B0",x"D7",x"B0",x"A4",x"80",x"27", -- 0xAC78
    x"E8",x"E6",x"42",x"E7",x"62",x"C6",x"F8",x"CB", -- 0xAC80
    x"08",x"44",x"24",x"FB",x"EB",x"E4",x"C1",x"1A", -- 0xAC88
    x"22",x"1D",x"0D",x"70",x"27",x"04",x"8D",x"44", -- 0xAC90
    x"26",x"02",x"CB",x"40",x"E7",x"E4",x"8D",x"AB", -- 0xAC98
    x"A6",x"62",x"8D",x"46",x"A1",x"61",x"26",x"03", -- 0xACA0
    x"E6",x"E4",x"8C",x"6F",x"E4",x"35",x"92",x"8E", -- 0xACA8
    x"CC",x"DE",x"C1",x"21",x"25",x"16",x"8E",x"CC", -- 0xACB0
    x"C0",x"C1",x"30",x"24",x"0F",x"8D",x"24",x"C1", -- 0xACB8
    x"2B",x"23",x"02",x"88",x"40",x"4D",x"26",x"D4", -- 0xACC0
    x"CB",x"10",x"20",x"D0",x"58",x"0D",x"70",x"27", -- 0xACC8
    x"02",x"CB",x"12",x"8D",x"0E",x"27",x"01",x"5C", -- 0xACD0
    x"E6",x"85",x"20",x"C0",x"86",x"EF",x"8D",x"24", -- 0xACD8
    x"84",x"08",x"39",x"86",x"7F",x"8D",x"1D",x"84", -- 0xACE0
    x"40",x"39",x"A7",x"42",x"8D",x"18",x"6D",x"42", -- 0xACE8
    x"2B",x"03",x"84",x"3F",x"39",x"0D",x"70",x"27", -- 0xACF0
    x"08",x"E6",x"42",x"C1",x"EF",x"26",x"02",x"84", -- 0xACF8
    x"77",x"1A",x"01",x"39",x"A7",x"42",x"0D",x"70", -- 0xAD00
    x"27",x"04",x"13",x"96",x"6A",x"8C",x"A6",x"C4", -- 0xAD08
    x"43",x"84",x"7F",x"39",x"0B",x"1B",x"0A",x"1A", -- 0xAD10
    x"08",x"18",x"09",x"19",x"20",x"20",x"30",x"5F", -- 0xAD18
    x"0D",x"1D",x"0C",x"1C",x"03",x"13",x"5E",x"5C", -- 0xAD20
    x"00",x"00",x"08",x"5B",x"09",x"5D",x"20",x"20", -- 0xAD28
    x"30",x"5F",x"0D",x"0D",x"1B",x"80",x"FF",x"8F", -- 0xAD30
    x"20",x"3F",x"54",x"50",x"4D",x"4F",x"52",x"50", -- 0xAD38
    x"4F",x"56",x"45",x"52",x"4C",x"41",x"50",x"3F", -- 0xAD40
    x"8D",x"02",x"1F",x"98",x"E6",x"01",x"54",x"54", -- 0xAD48
    x"54",x"54",x"EA",x"81",x"39",x"6F",x"84",x"8C", -- 0xAD50
    x"6C",x"84",x"A3",x"63",x"24",x"FA",x"E3",x"63", -- 0xAD58
    x"39",x"A6",x"49",x"8B",x"0F",x"D6",x"66",x"3D", -- 0xAD60
    x"97",x"1C",x"30",x"41",x"8D",x"DA",x"DD",x"18", -- 0xAD68
    x"8D",x"D6",x"DD",x"1A",x"DC",x"18",x"26",x"04", -- 0xAD70
    x"DC",x"1A",x"DD",x"18",x"D3",x"18",x"24",x"04", -- 0xAD78
    x"98",x"1A",x"D8",x"1B",x"DD",x"18",x"84",x"80", -- 0xAD80
    x"27",x"02",x"96",x"1C",x"A7",x"9F",x"00",x"16", -- 0xAD88
    x"0C",x"17",x"26",x"E0",x"7E",x"CE",x"5A",x"34", -- 0xAD90
    x"14",x"8E",x"00",x"6B",x"1F",x"89",x"4F",x"8D", -- 0xAD98
    x"B4",x"1F",x"98",x"E6",x"E4",x"30",x"01",x"8D", -- 0xADA0
    x"AC",x"35",x"14",x"DC",x"6B",x"39",x"BD",x"DA", -- 0xADA8
    x"E4",x"8E",x"CE",x"E2",x"CE",x"08",x"00",x"BD", -- 0xADB0
    x"D4",x"AA",x"35",x"20",x"C6",x"80",x"30",x"85", -- 0xADB8
    x"A6",x"80",x"40",x"A7",x"C0",x"5A",x"26",x"F8", -- 0xADC0
    x"0F",x"56",x"10",x"8E",x"0F",x"00",x"86",x"0A", -- 0xADC8
    x"97",x"16",x"CC",x"0A",x"04",x"97",x"6C",x"A6", -- 0xADD0
    x"A0",x"A1",x"A8",x"31",x"34",x"01",x"E4",x"E0", -- 0xADD8
    x"A7",x"A8",x"31",x"0A",x"6C",x"26",x"F0",x"5D", -- 0xADE0
    x"26",x"70",x"0F",x"17",x"33",x"36",x"6D",x"C4", -- 0xADE8
    x"10",x"27",x"FF",x"6D",x"86",x"08",x"9E",x"8A", -- 0xADF0
    x"9F",x"14",x"E6",x"C6",x"3A",x"4A",x"26",x"FA", -- 0xADF8
    x"86",x"08",x"34",x"02",x"5F",x"A6",x"C6",x"27", -- 0xAE00
    x"07",x"8D",x"8C",x"4A",x"2B",x"02",x"C6",x"FF", -- 0xAE08
    x"35",x"02",x"E7",x"C6",x"4A",x"26",x"EB",x"8D", -- 0xAE10
    x"6A",x"4D",x"2A",x"02",x"8D",x"57",x"10",x"93", -- 0xAE18
    x"14",x"25",x"02",x"DD",x"14",x"0C",x"17",x"2A", -- 0xAE20
    x"EE",x"DC",x"14",x"8D",x"4F",x"34",x"06",x"AE", -- 0xAE28
    x"E1",x"27",x"06",x"96",x"67",x"5F",x"BD",x"CD", -- 0xAE30
    x"97",x"D7",x"14",x"0F",x"17",x"8D",x"44",x"D6", -- 0xAE38
    x"14",x"8D",x"2D",x"8D",x"37",x"1F",x"98",x"E6", -- 0xAE40
    x"49",x"CB",x"0F",x"8D",x"23",x"9B",x"67",x"2A", -- 0xAE48
    x"01",x"4F",x"A7",x"9F",x"00",x"16",x"0C",x"17", -- 0xAE50
    x"26",x"E3",x"96",x"16",x"4C",x"81",x"0F",x"10", -- 0xAE58
    x"25",x"FF",x"6D",x"0D",x"5A",x"26",x"48",x"0D", -- 0xAE60
    x"59",x"27",x"41",x"BD",x"C9",x"0D",x"20",x"3F", -- 0xAE68
    x"4D",x"2A",x"6C",x"40",x"3D",x"53",x"43",x"C9", -- 0xAE70
    x"00",x"89",x"00",x"39",x"8D",x"00",x"8D",x"00", -- 0xAE78
    x"47",x"56",x"39",x"6F",x"E2",x"6F",x"E2",x"86", -- 0xAE80
    x"08",x"34",x"02",x"E6",x"C6",x"27",x"16",x"34", -- 0xAE88
    x"04",x"5F",x"DB",x"17",x"4A",x"26",x"FB",x"8E", -- 0xAE90
    x"08",x"00",x"3A",x"A6",x"84",x"35",x"04",x"8D", -- 0xAE98
    x"CF",x"E3",x"61",x"ED",x"61",x"35",x"02",x"4A", -- 0xAEA0
    x"26",x"DF",x"35",x"86",x"BD",x"C9",x"2F",x"0F", -- 0xAEA8
    x"5D",x"0F",x"59",x"10",x"CE",x"00",x"F8",x"1A", -- 0xAEB0
    x"FF",x"1F",x"AB",x"0F",x"D8",x"0F",x"D6",x"0F", -- 0xAEB8
    x"C6",x"CC",x"35",x"3C",x"97",x"01",x"D7",x"03", -- 0xAEC0
    x"4A",x"97",x"21",x"D7",x"23",x"0D",x"02",x"0F", -- 0xAEC8
    x"22",x"CC",x"00",x"03",x"DA",x"7F",x"D7",x"7F", -- 0xAED0
    x"0F",x"40",x"1F",x"8B",x"0F",x"A0",x"39",x"3D", -- 0xAED8
    x"39",x"80",x"00",x"01",x"02",x"03",x"04",x"05", -- 0xAEE0
    x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D", -- 0xAEE8
    x"0E",x"0F",x"10",x"11",x"12",x"13",x"14",x"15", -- 0xAEF0
    x"16",x"17",x"18",x"18",x"19",x"1A",x"1B",x"1C", -- 0xAEF8
    x"1C",x"1D",x"1E",x"1F",x"1F",x"20",x"21",x"21", -- 0xAF00
    x"22",x"23",x"23",x"24",x"24",x"25",x"25",x"26", -- 0xAF08
    x"26",x"27",x"27",x"27",x"28",x"28",x"29",x"29", -- 0xAF10
    x"29",x"29",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A", -- 0xAF18
    x"2A",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A", -- 0xAF20
    x"2A",x"2A",x"2A",x"29",x"29",x"29",x"29",x"28", -- 0xAF28
    x"28",x"27",x"27",x"27",x"26",x"26",x"25",x"25", -- 0xAF30
    x"24",x"24",x"23",x"23",x"22",x"21",x"21",x"20", -- 0xAF38
    x"1F",x"1F",x"1E",x"1D",x"1C",x"1C",x"1B",x"1A", -- 0xAF40
    x"19",x"18",x"18",x"17",x"16",x"15",x"14",x"13", -- 0xAF48
    x"12",x"11",x"10",x"0F",x"0E",x"0D",x"0C",x"0B", -- 0xAF50
    x"0A",x"09",x"08",x"07",x"06",x"05",x"04",x"03", -- 0xAF58
    x"02",x"01",x"00",x"02",x"03",x"05",x"06",x"08", -- 0xAF60
    x"09",x"0B",x"0C",x"0E",x"0F",x"11",x"12",x"14", -- 0xAF68
    x"15",x"17",x"18",x"1A",x"1B",x"1D",x"1E",x"1F", -- 0xAF70
    x"21",x"22",x"23",x"25",x"26",x"27",x"28",x"29", -- 0xAF78
    x"2B",x"2C",x"2D",x"2E",x"2F",x"30",x"31",x"32", -- 0xAF80
    x"33",x"34",x"35",x"36",x"36",x"37",x"38",x"39", -- 0xAF88
    x"39",x"3A",x"3B",x"3B",x"3C",x"3C",x"3D",x"3D", -- 0xAF90
    x"3E",x"3E",x"3E",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0xAF98
    x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0xAFA0
    x"3F",x"3F",x"3E",x"3E",x"3E",x"3D",x"3D",x"3C", -- 0xAFA8
    x"3C",x"3B",x"3B",x"3A",x"39",x"39",x"38",x"37", -- 0xAFB0
    x"36",x"36",x"35",x"34",x"33",x"32",x"31",x"30", -- 0xAFB8
    x"2F",x"2E",x"2D",x"2C",x"2B",x"29",x"28",x"27", -- 0xAFC0
    x"26",x"25",x"23",x"22",x"21",x"1F",x"1E",x"1D", -- 0xAFC8
    x"1B",x"1A",x"18",x"17",x"15",x"14",x"12",x"11", -- 0xAFD0
    x"0F",x"0E",x"0C",x"0B",x"09",x"08",x"06",x"05", -- 0xAFD8
    x"03",x"02",x"71",x"29",x"72",x"12",x"73",x"B4", -- 0xAFE0
    x"76",x"57",x"FF",x"01",x"E0",x"F0",x"A0",x"50", -- 0xAFE8
    x"40",x"40",x"00",x"00",x"E0",x"01",x"40",x"80", -- 0xAFF0
    x"F0",x"80",x"F0",x"20",x"00",x"00",x"F0",x"01", -- 0xAFF8
    x"E0",x"00",x"50",x"00",x"F0",x"00",x"00",x"00", -- 0xB000
    x"A0",x"01",x"F0",x"40",x"00",x"80",x"00",x"00", -- 0xB008
    x"00",x"00",x"B0",x"01",x"40",x"F0",x"20",x"80", -- 0xB010
    x"10",x"40",x"00",x"00",x"D0",x"29",x"2A",x"2C", -- 0xB018
    x"68",x"0F",x"A9",x"39",x"7E",x"D2",x"06",x"0F", -- 0xB020
    x"8E",x"CC",x"01",x"20",x"97",x"A1",x"A6",x"A5", -- 0xB028
    x"4C",x"26",x"1D",x"E7",x"C4",x"33",x"A5",x"86", -- 0xB030
    x"C0",x"A7",x"C4",x"34",x"04",x"1F",x"98",x"44", -- 0xB038
    x"81",x"11",x"25",x"01",x"4C",x"C4",x"01",x"27", -- 0xB040
    x"02",x"C6",x"09",x"5C",x"DD",x"A3",x"35",x"84", -- 0xB048
    x"DB",x"A1",x"2B",x"D0",x"C1",x"44",x"26",x"D6", -- 0xB050
    x"00",x"A1",x"C6",x"1F",x"20",x"D0",x"0C",x"5B", -- 0xB058
    x"BD",x"D2",x"FB",x"BD",x"D3",x"89",x"BD",x"D3", -- 0xB060
    x"70",x"25",x"B9",x"A6",x"84",x"27",x"03",x"4C", -- 0xB068
    x"26",x"F4",x"CE",x"00",x"0D",x"8D",x"B0",x"DC", -- 0xB070
    x"5E",x"DD",x"7E",x"86",x"20",x"97",x"9F",x"86", -- 0xB078
    x"08",x"91",x"8E",x"24",x"02",x"8D",x"A0",x"BD", -- 0xB080
    x"D3",x"AB",x"0C",x"7E",x"0C",x"A4",x"0C",x"8E", -- 0xB088
    x"0A",x"0E",x"2A",x"EB",x"0C",x"0E",x"96",x"8E", -- 0xB090
    x"8A",x"C0",x"A7",x"C4",x"9E",x"8A",x"DE",x"8C", -- 0xB098
    x"C6",x"10",x"BD",x"D4",x"B1",x"7E",x"D3",x"22", -- 0xB0A0
    x"9E",x"5E",x"8D",x"45",x"10",x"2B",x"FB",x"01", -- 0xB0A8
    x"DC",x"74",x"93",x"5E",x"DD",x"0E",x"0D",x"A9", -- 0xB0B0
    x"26",x"A4",x"AD",x"9F",x"A0",x"0C",x"8D",x"2D", -- 0xB0B8
    x"CC",x"50",x"FF",x"4A",x"26",x"FD",x"4C",x"DD", -- 0xB0C0
    x"7C",x"9E",x"12",x"CE",x"08",x"02",x"DF",x"7E", -- 0xB0C8
    x"BD",x"D4",x"B1",x"9F",x"12",x"CC",x"FF",x"01", -- 0xB0D0
    x"D3",x"0E",x"DD",x"0E",x"2A",x"E0",x"C3",x"00", -- 0xB0D8
    x"FF",x"D7",x"7D",x"27",x"03",x"4D",x"2A",x"D6", -- 0xB0E0
    x"CC",x"FF",x"00",x"DD",x"7C",x"6E",x"9F",x"A0", -- 0xB0E8
    x"08",x"9F",x"12",x"BD",x"C9",x"08",x"BD",x"D7", -- 0xB0F0
    x"0D",x"DF",x"64",x"9E",x"8A",x"9F",x"A1",x"CC", -- 0xB0F8
    x"00",x"0F",x"DD",x"7C",x"86",x"20",x"A7",x"80", -- 0xB100
    x"5A",x"2A",x"FB",x"86",x"01",x"DD",x"0B",x"0F", -- 0xB108
    x"0D",x"9E",x"8A",x"0D",x"A9",x"26",x"02",x"30", -- 0xB110
    x"03",x"9F",x"7E",x"E7",x"84",x"C6",x"08",x"A6", -- 0xB118
    x"C0",x"2B",x"31",x"81",x"60",x"27",x"2D",x"81", -- 0xB120
    x"7A",x"27",x"1D",x"81",x"6F",x"27",x"11",x"85", -- 0xB128
    x"20",x"27",x"02",x"84",x"BF",x"A7",x"80",x"81", -- 0xB130
    x"2A",x"26",x"02",x"97",x"A1",x"5A",x"26",x"DF", -- 0xB138
    x"A6",x"C0",x"2B",x"10",x"81",x"7A",x"26",x"F8", -- 0xB140
    x"A6",x"C0",x"80",x"70",x"81",x"04",x"97",x"A2", -- 0xB148
    x"10",x"24",x"00",x"B2",x"96",x"03",x"9A",x"00", -- 0xB150
    x"2B",x"06",x"0D",x"A1",x"26",x"02",x"0F",x"A7", -- 0xB158
    x"4D",x"39",x"0D",x"A9",x"10",x"26",x"FA",x"9A", -- 0xB160
    x"21",x"CC",x"DC",x"8A",x"9E",x"74",x"20",x"04", -- 0xB168
    x"9E",x"5E",x"4F",x"5C",x"DD",x"6B",x"BD",x"D0", -- 0xB170
    x"F1",x"10",x"2B",x"FA",x"34",x"8E",x"08",x"02", -- 0xB178
    x"9F",x"7E",x"0D",x"6B",x"27",x"03",x"BD",x"C9", -- 0xB180
    x"2B",x"0D",x"A9",x"10",x"26",x"00",x"C5",x"8E", -- 0xB188
    x"04",x"20",x"CC",x"0F",x"13",x"E7",x"80",x"BD", -- 0xB190
    x"C9",x"1B",x"AD",x"9F",x"A0",x"04",x"8D",x"6A", -- 0xB198
    x"0D",x"7C",x"2B",x"E5",x"26",x"F4",x"CE",x"04", -- 0xB1A0
    x"22",x"BD",x"D3",x"08",x"30",x"18",x"CE",x"00", -- 0xB1A8
    x"03",x"C6",x"08",x"A6",x"C0",x"81",x"2A",x"27", -- 0xB1B0
    x"07",x"A1",x"80",x"26",x"DD",x"5A",x"26",x"F3", -- 0xB1B8
    x"3A",x"EE",x"84",x"11",x"93",x"0B",x"26",x"D2", -- 0xB1C0
    x"0D",x"81",x"26",x"3A",x"EE",x"03",x"DF",x"0E", -- 0xB1C8
    x"DC",x"12",x"93",x"0E",x"25",x"43",x"10",x"83", -- 0xB1D0
    x"10",x"64",x"23",x"3D",x"1F",x"03",x"0D",x"6C", -- 0xB1D8
    x"27",x"02",x"DF",x"5E",x"11",x"93",x"5E",x"26", -- 0xB1E0
    x"1D",x"86",x"46",x"B7",x"04",x"20",x"DF",x"12", -- 0xB1E8
    x"8D",x"18",x"4D",x"26",x"11",x"0D",x"7C",x"27", -- 0xB1F0
    x"0D",x"2B",x"45",x"DE",x"12",x"D6",x"7D",x"27", -- 0xB1F8
    x"ED",x"BD",x"D4",x"95",x"27",x"E8",x"86",x"77", -- 0xB200
    x"20",x"17",x"B6",x"04",x"20",x"88",x"40",x"B7", -- 0xB208
    x"04",x"20",x"AD",x"9F",x"A0",x"06",x"9E",x"7E", -- 0xB210
    x"39",x"86",x"71",x"0D",x"59",x"27",x"02",x"0F", -- 0xB218
    x"56",x"B7",x"04",x"3E",x"CC",x"45",x"52",x"F7", -- 0xB220
    x"04",x"3C",x"FD",x"04",x"3A",x"0D",x"56",x"27", -- 0xB228
    x"05",x"30",x"5F",x"BD",x"C8",x"E3",x"0D",x"59", -- 0xB230
    x"27",x"03",x"BD",x"C9",x"0D",x"7E",x"DD",x"A4", -- 0xB238
    x"9E",x"5E",x"86",x"8F",x"B7",x"04",x"20",x"7E", -- 0xB240
    x"C9",x"2D",x"0D",x"58",x"27",x"B8",x"0D",x"A7", -- 0xB248
    x"27",x"B4",x"0F",x"A7",x"8D",x"6B",x"25",x"F2", -- 0xB250
    x"C6",x"03",x"8D",x"60",x"30",x"10",x"CE",x"04", -- 0xB258
    x"22",x"BD",x"D3",x"08",x"1F",x"31",x"BD",x"C9", -- 0xB260
    x"19",x"8E",x"0F",x"64",x"9F",x"02",x"D6",x"0D", -- 0xB268
    x"2B",x"29",x"BD",x"D0",x"3B",x"86",x"09",x"E6", -- 0xB270
    x"A5",x"D7",x"0D",x"2A",x"06",x"1F",x"98",x"84", -- 0xB278
    x"0F",x"27",x"83",x"97",x"8E",x"DC",x"02",x"4C", -- 0xB280
    x"10",x"93",x"12",x"24",x"8C",x"5F",x"8D",x"28", -- 0xB288
    x"BD",x"D3",x"AB",x"0C",x"A4",x"0A",x"8E",x"26", -- 0xB290
    x"EC",x"20",x"D3",x"DC",x"0E",x"27",x"02",x"8D", -- 0xB298
    x"17",x"8E",x"10",x"64",x"9F",x"5E",x"9E",x"12", -- 0xB2A0
    x"8D",x"02",x"20",x"96",x"A6",x"C2",x"8A",x"40", -- 0xB2A8
    x"A7",x"82",x"11",x"93",x"5E",x"22",x"F5",x"39", -- 0xB2B0
    x"9E",x"7E",x"DE",x"02",x"8D",x"37",x"DF",x"02", -- 0xB2B8
    x"39",x"53",x"06",x"5B",x"BD",x"D3",x"8B",x"BD", -- 0xB2C0
    x"D3",x"70",x"25",x"47",x"6D",x"84",x"2F",x"F7", -- 0xB2C8
    x"CE",x"00",x"08",x"30",x"08",x"C6",x"05",x"BD", -- 0xB2D0
    x"D4",x"99",x"26",x"EB",x"DE",x"8A",x"30",x"13", -- 0xB2D8
    x"C6",x"0D",x"BD",x"D4",x"99",x"27",x"2C",x"0D", -- 0xB2E0
    x"5B",x"2A",x"DC",x"81",x"2A",x"26",x"D8",x"97", -- 0xB2E8
    x"A7",x"30",x"1F",x"33",x"5F",x"7E",x"D4",x"B1", -- 0xB2F0
    x"BD",x"D0",x"F1",x"0F",x"A7",x"8D",x"C5",x"24", -- 0xB2F8
    x"13",x"0D",x"5B",x"26",x"0E",x"7E",x"D2",x"06", -- 0xB300
    x"C6",x"08",x"A6",x"80",x"8A",x"40",x"A7",x"C0", -- 0xB308
    x"5A",x"26",x"F7",x"39",x"A6",x"84",x"E6",x"A6", -- 0xB310
    x"6F",x"A6",x"6A",x"A6",x"E7",x"84",x"2A",x"F4", -- 0xB318
    x"6F",x"13",x"8D",x"78",x"86",x"20",x"8E",x"09", -- 0xB320
    x"00",x"C6",x"02",x"20",x"76",x"5C",x"D7",x"A9", -- 0xB328
    x"0F",x"A2",x"BD",x"D7",x"0D",x"2B",x"03",x"BD", -- 0xB330
    x"D0",x"F1",x"8D",x"4D",x"8E",x"04",x"40",x"1F", -- 0xB338
    x"13",x"86",x"0E",x"BD",x"C9",x"1B",x"8D",x"28", -- 0xB340
    x"25",x"C9",x"A6",x"84",x"2F",x"F8",x"A6",x"08", -- 0xB348
    x"E6",x"0B",x"E4",x"0C",x"10",x"83",x"20",x"01", -- 0xB350
    x"26",x"EC",x"8D",x"AC",x"1F",x"30",x"C5",x"1F", -- 0xB358
    x"27",x"02",x"33",x"44",x"11",x"93",x"AD",x"25", -- 0xB360
    x"DD",x"BD",x"CC",x"5B",x"27",x"FB",x"20",x"CC", -- 0xB368
    x"9E",x"8C",x"30",x"88",x"20",x"8C",x"09",x"00", -- 0xB370
    x"25",x"0B",x"0C",x"A6",x"D6",x"A6",x"C1",x"0C", -- 0xB378
    x"24",x"14",x"4F",x"8D",x"19",x"4F",x"9F",x"8C", -- 0xB380
    x"39",x"0F",x"A7",x"4F",x"8D",x"98",x"1F",x"12", -- 0xB388
    x"0D",x"A7",x"26",x"0A",x"9F",x"8C",x"86",x"02", -- 0xB390
    x"97",x"A6",x"43",x"39",x"86",x"20",x"8E",x"08", -- 0xB398
    x"00",x"D6",x"A6",x"97",x"9F",x"86",x"11",x"DD", -- 0xB3A0
    x"A3",x"9F",x"7E",x"34",x"74",x"CE",x"FF",x"40", -- 0xB3A8
    x"C6",x"04",x"D7",x"6B",x"DC",x"A2",x"8E",x"D0", -- 0xB3B0
    x"1D",x"A6",x"86",x"C1",x"16",x"25",x"02",x"8A", -- 0xB3B8
    x"10",x"A7",x"C4",x"0D",x"A0",x"26",x"04",x"8D", -- 0xB3C0
    x"3F",x"8D",x"3D",x"97",x"A0",x"8D",x"29",x"26", -- 0xB3C8
    x"04",x"0F",x"A5",x"8D",x"49",x"96",x"A5",x"27", -- 0xB3D0
    x"0C",x"0A",x"6B",x"10",x"27",x"FE",x"27",x"8D", -- 0xB3D8
    x"06",x"26",x"F2",x"20",x"CF",x"35",x"F4",x"8E", -- 0xB3E0
    x"00",x"FC",x"D6",x"A2",x"6F",x"85",x"86",x"03", -- 0xB3E8
    x"8D",x"04",x"84",x"10",x"20",x"25",x"8D",x"15", -- 0xB3F0
    x"9E",x"8A",x"30",x"1F",x"27",x"15",x"A6",x"48", -- 0xB3F8
    x"85",x"01",x"26",x"F6",x"39",x"8E",x"23",x"45", -- 0xB400
    x"30",x"1F",x"26",x"FC",x"39",x"A7",x"48",x"34", -- 0xB408
    x"06",x"35",x"86",x"86",x"D0",x"8D",x"F6",x"A6", -- 0xB410
    x"48",x"8A",x"80",x"97",x"A5",x"39",x"8E",x"00", -- 0xB418
    x"FC",x"D6",x"A2",x"A6",x"85",x"A7",x"49",x"91", -- 0xB420
    x"A3",x"27",x"12",x"96",x"A3",x"A7",x"4B",x"A7", -- 0xB428
    x"85",x"86",x"17",x"8D",x"C1",x"26",x"E6",x"8D", -- 0xB430
    x"CC",x"84",x"18",x"26",x"DE",x"D6",x"A4",x"E7", -- 0xB438
    x"4A",x"9E",x"7E",x"10",x"9E",x"8A",x"6D",x"48", -- 0xB440
    x"CC",x"80",x"80",x"D3",x"9F",x"81",x"A0",x"8D", -- 0xB448
    x"BC",x"86",x"02",x"97",x"A8",x"25",x"14",x"A5", -- 0xB450
    x"48",x"26",x"08",x"31",x"3F",x"26",x"F8",x"0F", -- 0xB458
    x"A8",x"20",x"B0",x"A6",x"80",x"A7",x"4B",x"E7", -- 0xB460
    x"C4",x"20",x"F8",x"A5",x"48",x"26",x"06",x"31", -- 0xB468
    x"3F",x"26",x"F8",x"20",x"EA",x"A6",x"4B",x"A7", -- 0xB470
    x"80",x"E7",x"C4",x"20",x"F8",x"7D",x"00",x"A8", -- 0xB478
    x"26",x"01",x"3B",x"32",x"6C",x"0F",x"A8",x"A6", -- 0xB480
    x"48",x"84",x"7C",x"20",x"8E",x"32",x"62",x"4F", -- 0xB488
    x"8D",x"4A",x"7E",x"CB",x"E6",x"0D",x"6C",x"26", -- 0xB490
    x"18",x"A6",x"C0",x"A1",x"80",x"26",x"03",x"5A", -- 0xB498
    x"26",x"F7",x"39",x"6D",x"C0",x"2A",x"FC",x"33", -- 0xB4A0
    x"5F",x"39",x"E6",x"1F",x"0D",x"AA",x"26",x"01", -- 0xB4A8
    x"3A",x"A6",x"80",x"A7",x"C0",x"5A",x"26",x"F9", -- 0xB4B0
    x"39",x"DE",x"5E",x"8D",x"E6",x"A6",x"C0",x"84", -- 0xB4B8
    x"7F",x"27",x"12",x"81",x"6F",x"27",x"F4",x"81", -- 0xB4C0
    x"56",x"26",x"F2",x"A6",x"C4",x"84",x"7F",x"81", -- 0xB4C8
    x"75",x"26",x"EA",x"80",x"74",x"97",x"AA",x"4F", -- 0xB4D0
    x"0F",x"78",x"0A",x"78",x"DD",x"76",x"0C",x"56", -- 0xB4D8
    x"8E",x"D5",x"22",x"CE",x"00",x"66",x"8D",x"C2", -- 0xB4E0
    x"8E",x"CF",x"EB",x"CE",x"0F",x"00",x"C6",x"32", -- 0xB4E8
    x"96",x"AA",x"91",x"AB",x"27",x"03",x"58",x"97", -- 0xB4F0
    x"AB",x"8D",x"B6",x"BD",x"DC",x"88",x"1E",x"31", -- 0xB4F8
    x"C6",x"39",x"BD",x"C9",x"F6",x"CE",x"D5",x"2A", -- 0xB500
    x"1E",x"13",x"C6",x"0A",x"8D",x"A3",x"8E",x"0F", -- 0xB508
    x"64",x"9F",x"51",x"AF",x"42",x"30",x"0C",x"9F", -- 0xB510
    x"7A",x"AF",x"C4",x"DE",x"5E",x"8D",x"24",x"20", -- 0xB518
    x"FC",x"04",x"55",x"2A",x"0A",x"05",x"7F",x"40", -- 0xB520
    x"06",x"04",x"00",x"00",x"00",x"0D",x"0D",x"0D", -- 0xB528
    x"0D",x"0D",x"02",x"60",x"48",x"60",x"49",x"18", -- 0xB530
    x"51",x"30",x"53",x"0C",x"54",x"06",x"57",x"C0", -- 0xB538
    x"58",x"03",x"FF",x"8D",x"60",x"4D",x"10",x"27", -- 0xB540
    x"F8",x"64",x"8E",x"D6",x"69",x"BD",x"CB",x"D1", -- 0xB548
    x"0D",x"53",x"26",x"EF",x"8E",x"D5",x"34",x"BD", -- 0xB550
    x"D6",x"50",x"25",x"2E",x"1F",x"89",x"D7",x"0E", -- 0xB558
    x"8D",x"43",x"81",x"7A",x"26",x"10",x"58",x"25", -- 0xB560
    x"17",x"4F",x"C0",x"03",x"4C",x"24",x"FB",x"4A", -- 0xB568
    x"1F",x"89",x"D7",x"0E",x"8D",x"2F",x"81",x"6E", -- 0xB570
    x"26",x"0B",x"04",x"0E",x"DB",x"0E",x"24",x"F4", -- 0xB578
    x"86",x"76",x"7E",x"D2",x"21",x"D7",x"0E",x"33", -- 0xB580
    x"5F",x"39",x"D6",x"12",x"BD",x"D6",x"B4",x"D7", -- 0xB588
    x"6C",x"8D",x"5E",x"8D",x"5C",x"C8",x"10",x"34", -- 0xB590
    x"04",x"CA",x"70",x"E1",x"E4",x"35",x"04",x"26", -- 0xB598
    x"20",x"D6",x"6C",x"20",x"1C",x"DF",x"62",x"A6", -- 0xB5A0
    x"C0",x"2A",x"10",x"33",x"5F",x"DF",x"60",x"11", -- 0xB5A8
    x"93",x"76",x"26",x"03",x"BD",x"DA",x"11",x"A6", -- 0xB5B0
    x"C0",x"84",x"7F",x"39",x"32",x"62",x"8C",x"C6", -- 0xB5B8
    x"70",x"86",x"FF",x"97",x"6C",x"9E",x"8A",x"96", -- 0xB5C0
    x"10",x"31",x"86",x"AE",x"A4",x"D7",x"6B",x"A6", -- 0xB5C8
    x"1F",x"91",x"6B",x"27",x"0E",x"84",x"8F",x"91", -- 0xB5D0
    x"6B",x"26",x"20",x"86",x"60",x"A4",x"1F",x"81", -- 0xB5D8
    x"60",x"27",x"18",x"A6",x"1E",x"9B",x"0E",x"25", -- 0xB5E0
    x"12",x"81",x"FF",x"27",x"0E",x"A7",x"1E",x"20", -- 0xB5E8
    x"14",x"8E",x"D6",x"59",x"8D",x"50",x"25",x"C4", -- 0xB5F0
    x"EA",x"1F",x"39",x"96",x"0E",x"A7",x"80",x"A6", -- 0xB5F8
    x"84",x"97",x"6C",x"E7",x"80",x"34",x"10",x"8E", -- 0xB600
    x"D6",x"60",x"8D",x"3A",x"35",x"10",x"25",x"2B", -- 0xB608
    x"44",x"24",x"08",x"1F",x"89",x"96",x"0E",x"44", -- 0xB610
    x"5A",x"26",x"FC",x"1F",x"89",x"40",x"27",x"1B", -- 0xB618
    x"AB",x"1E",x"A7",x"1E",x"96",x"12",x"48",x"27", -- 0xB620
    x"06",x"A6",x"1E",x"E7",x"1E",x"1F",x"89",x"E7", -- 0xB628
    x"80",x"A6",x"84",x"C6",x"70",x"E7",x"80",x"94", -- 0xB630
    x"6C",x"97",x"6C",x"AF",x"A4",x"0C",x"6C",x"27", -- 0xB638
    x"B9",x"86",x"75",x"7E",x"D2",x"21",x"BD",x"D5", -- 0xB640
    x"A5",x"8D",x"05",x"24",x"0B",x"33",x"5F",x"39", -- 0xB648
    x"A1",x"81",x"25",x"04",x"26",x"FA",x"A6",x"1F", -- 0xB650
    x"39",x"63",x"20",x"65",x"10",x"66",x"40",x"FF", -- 0xB658
    x"62",x"04",x"67",x"02",x"6C",x"03",x"7B",x"05", -- 0xB660
    x"FF",x"40",x"D6",x"DB",x"4A",x"D7",x"D4",x"4B", -- 0xB668
    x"D7",x"2B",x"4D",x"D6",x"F4",x"4E",x"D7",x"87", -- 0xB670
    x"4F",x"D7",x"9D",x"50",x"D8",x"3D",x"52",x"D8", -- 0xB678
    x"2D",x"55",x"D6",x"E2",x"56",x"D7",x"C7",x"59", -- 0xB680
    x"D7",x"59",x"5A",x"D7",x"B3",x"5F",x"D6",x"D8", -- 0xB688
    x"60",x"D7",x"86",x"64",x"D5",x"BF",x"68",x"D7", -- 0xB690
    x"71",x"69",x"D7",x"78",x"6A",x"D6",x"DE",x"6F", -- 0xB698
    x"D4",x"A3",x"7C",x"D7",x"AE",x"7D",x"D7",x"BF", -- 0xB6A0
    x"7E",x"D7",x"98",x"FF",x"6B",x"00",x"6D",x"80", -- 0xB6A8
    x"FF",x"BD",x"D5",x"A5",x"34",x"04",x"8E",x"D6", -- 0xB6B0
    x"AC",x"8D",x"95",x"25",x"05",x"A7",x"E4",x"BD", -- 0xB6B8
    x"D5",x"A5",x"81",x"47",x"26",x"04",x"6D",x"E4", -- 0xB6C0
    x"2A",x"0C",x"BD",x"D7",x"FB",x"4D",x"26",x"02", -- 0xB6C8
    x"8A",x"80",x"AA",x"E4",x"A7",x"E4",x"35",x"84", -- 0xB6D0
    x"86",x"E0",x"8C",x"86",x"80",x"21",x"4F",x"97", -- 0xB6D8
    x"12",x"39",x"C6",x"80",x"8D",x"CB",x"8E",x"00", -- 0xB6E0
    x"0D",x"96",x"10",x"5D",x"2A",x"03",x"C8",x"7F", -- 0xB6E8
    x"5C",x"E7",x"86",x"39",x"34",x"40",x"BD",x"DB", -- 0xB6F0
    x"25",x"0D",x"17",x"26",x"0B",x"8E",x"00",x"19", -- 0xB6F8
    x"CE",x"00",x"20",x"C6",x"23",x"BD",x"D4",x"B1", -- 0xB700
    x"35",x"40",x"0F",x"17",x"8C",x"33",x"21",x"A6", -- 0xB708
    x"C0",x"2B",x"0A",x"81",x"60",x"26",x"F8",x"A6", -- 0xB710
    x"C0",x"81",x"60",x"27",x"FA",x"6D",x"C2",x"39", -- 0xB718
    x"48",x"01",x"49",x"04",x"51",x"02",x"53",x"08", -- 0xB720
    x"54",x"10",x"FF",x"8E",x"00",x"19",x"C6",x"07", -- 0xB728
    x"BD",x"C9",x"F6",x"BD",x"D5",x"A5",x"80",x"70", -- 0xB730
    x"81",x"08",x"24",x"57",x"1F",x"89",x"BD",x"D5", -- 0xB738
    x"A5",x"81",x"66",x"27",x"0D",x"30",x"19",x"81", -- 0xB740
    x"63",x"26",x"48",x"5A",x"2B",x"17",x"6C",x"80", -- 0xB748
    x"20",x"F9",x"5A",x"2B",x"10",x"6A",x"82",x"20", -- 0xB750
    x"F9",x"8D",x"0B",x"8B",x"0A",x"D6",x"10",x"54", -- 0xB758
    x"8E",x"00",x"46",x"A7",x"85",x"39",x"BD",x"D5", -- 0xB760
    x"A5",x"80",x"41",x"81",x"05",x"25",x"17",x"20", -- 0xB768
    x"22",x"DF",x"0A",x"86",x"FF",x"97",x"0C",x"39", -- 0xB770
    x"8D",x"7F",x"0D",x"0C",x"27",x"08",x"2A",x"02", -- 0xB778
    x"97",x"0C",x"0A",x"0C",x"DE",x"0A",x"39",x"8E", -- 0xB780
    x"D7",x"20",x"BD",x"D6",x"46",x"97",x"4B",x"24", -- 0xB788
    x"1C",x"33",x"41",x"86",x"73",x"7E",x"D2",x"21", -- 0xB790
    x"8D",x"5F",x"97",x"14",x"39",x"8D",x"5A",x"1F", -- 0xB798
    x"89",x"27",x"08",x"9A",x"16",x"84",x"01",x"DA", -- 0xB7A0
    x"17",x"C4",x"02",x"DD",x"16",x"39",x"8D",x"E8", -- 0xB7A8
    x"00",x"14",x"39",x"8D",x"44",x"91",x"68",x"24", -- 0xB7B0
    x"DA",x"C6",x"05",x"3D",x"D7",x"18",x"39",x"8D", -- 0xB7B8
    x"4B",x"44",x"27",x"CF",x"97",x"4C",x"39",x"BD", -- 0xB7C0
    x"D5",x"A5",x"80",x"71",x"81",x"05",x"24",x"C3", -- 0xB7C8
    x"48",x"97",x"10",x"39",x"8D",x"90",x"C6",x"0A", -- 0xB7D0
    x"3D",x"8E",x"0F",x"00",x"3A",x"BD",x"D5",x"A5", -- 0xB7D8
    x"80",x"52",x"81",x"02",x"24",x"E8",x"A7",x"80", -- 0xB7E0
    x"C6",x"09",x"8D",x"0D",x"48",x"48",x"48",x"48", -- 0xB7E8
    x"A7",x"80",x"5A",x"26",x"F5",x"39",x"1C",x"FB", -- 0xB7F0
    x"39",x"A6",x"C0",x"84",x"3F",x"80",x"30",x"81", -- 0xB7F8
    x"0A",x"25",x"08",x"8B",x"2F",x"81",x"06",x"24", -- 0xB800
    x"4D",x"8B",x"0A",x"39",x"BD",x"D5",x"A5",x"33", -- 0xB808
    x"5F",x"8D",x"E6",x"48",x"48",x"48",x"48",x"34", -- 0xB810
    x"02",x"8D",x"DE",x"AA",x"E0",x"39",x"8E",x"0F", -- 0xB818
    x"64",x"8C",x"AE",x"84",x"27",x"D0",x"9F",x"7C", -- 0xB820
    x"A1",x"02",x"26",x"F6",x"39",x"BD",x"DA",x"E4", -- 0xB828
    x"8D",x"DA",x"27",x"1F",x"8D",x"E8",x"26",x"1B", -- 0xB830
    x"AE",x"0A",x"9F",x"4D",x"39",x"BD",x"DA",x"E4", -- 0xB838
    x"BD",x"D5",x"A5",x"0F",x"45",x"81",x"60",x"27", -- 0xB840
    x"F3",x"8D",x"C4",x"97",x"45",x"27",x"ED",x"8D", -- 0xB848
    x"CD",x"26",x"E9",x"86",x"74",x"8C",x"86",x"72", -- 0xB850
    x"7E",x"D2",x"21",x"0F",x"56",x"0D",x"5D",x"26", -- 0xB858
    x"F2",x"BD",x"D7",x"0D",x"2B",x"03",x"8D",x"A9", -- 0xB860
    x"21",x"4F",x"8D",x"B2",x"26",x"E5",x"8E",x"DA", -- 0xB868
    x"7A",x"CE",x"08",x"9A",x"0D",x"5C",x"27",x"03", -- 0xB870
    x"33",x"C8",x"18",x"1F",x"32",x"BD",x"D4",x"AA", -- 0xB878
    x"EC",x"A8",x"16",x"44",x"56",x"ED",x"A3",x"10", -- 0xB880
    x"8C",x"08",x"22",x"26",x"F3",x"6F",x"A2",x"6F", -- 0xB888
    x"A2",x"EC",x"1E",x"0D",x"5C",x"27",x"02",x"47", -- 0xB890
    x"56",x"ED",x"A3",x"47",x"56",x"E3",x"A4",x"10", -- 0xB898
    x"8C",x"08",x"00",x"26",x"F4",x"CC",x"7F",x"EC", -- 0xB8A0
    x"ED",x"A4",x"CE",x"08",x"B4",x"8E",x"D8",x"E9", -- 0xB8A8
    x"BD",x"D4",x"AA",x"1F",x"31",x"CE",x"DA",x"AE", -- 0xB8B0
    x"96",x"AA",x"48",x"A6",x"C6",x"34",x"04",x"3D", -- 0xB8B8
    x"35",x"04",x"0D",x"5C",x"27",x"01",x"48",x"A7", -- 0xB8C0
    x"85",x"26",x"02",x"6C",x"85",x"5C",x"2A",x"E8", -- 0xB8C8
    x"10",x"8E",x"00",x"7C",x"CC",x"08",x"FB",x"F7", -- 0xB8D0
    x"FF",x"02",x"0D",x"5C",x"1F",x"8B",x"27",x"06", -- 0xB8D8
    x"7C",x"FF",x"D7",x"7C",x"FF",x"D9",x"0E",x"B4", -- 0xB8E0
    x"9C",x"20",x"61",x"86",x"00",x"A6",x"86",x"97", -- 0xB8E8
    x"B2",x"DC",x"20",x"C3",x"00",x"00",x"DD",x"BF", -- 0xB8F0
    x"97",x"EB",x"DC",x"20",x"C3",x"00",x"00",x"DD", -- 0xB8F8
    x"C8",x"97",x"EE",x"DC",x"20",x"C3",x"00",x"00", -- 0xB900
    x"DD",x"D1",x"97",x"F1",x"DC",x"20",x"C3",x"00", -- 0xB908
    x"00",x"DD",x"DA",x"97",x"F4",x"DC",x"20",x"C3", -- 0xB910
    x"00",x"00",x"DD",x"E3",x"97",x"F7",x"B6",x"0A", -- 0xB918
    x"00",x"BB",x"0A",x"00",x"F6",x"0A",x"00",x"FB", -- 0xB920
    x"0A",x"00",x"FB",x"0A",x"00",x"FD",x"FF",x"7A", -- 0xB928
    x"0A",x"B2",x"26",x"BD",x"0A",x"B3",x"26",x"08", -- 0xB930
    x"0A",x"B4",x"27",x"2E",x"96",x"B5",x"97",x"B3", -- 0xB938
    x"B6",x"FF",x"00",x"43",x"48",x"27",x"A4",x"2A", -- 0xB940
    x"A4",x"7E",x"DD",x"87",x"10",x"AE",x"A4",x"26", -- 0xB948
    x"03",x"7E",x"CE",x"B3",x"EC",x"23",x"97",x"EA", -- 0xB950
    x"D7",x"ED",x"EC",x"25",x"97",x"F0",x"D7",x"F3", -- 0xB958
    x"A6",x"27",x"97",x"F6",x"A6",x"29",x"97",x"B7", -- 0xB960
    x"EE",x"2A",x"37",x"06",x"97",x"B5",x"4C",x"27", -- 0xB968
    x"DB",x"D7",x"BD",x"37",x"06",x"97",x"C6",x"D7", -- 0xB970
    x"CF",x"37",x"06",x"97",x"D8",x"D7",x"E1",x"A6", -- 0xB978
    x"28",x"97",x"B4",x"20",x"B7",x"20",x"6E",x"86", -- 0xB980
    x"00",x"97",x"B3",x"B6",x"FF",x"00",x"43",x"48", -- 0xB988
    x"27",x"05",x"2A",x"05",x"7E",x"DD",x"87",x"86", -- 0xB990
    x"00",x"A6",x"86",x"97",x"B2",x"DC",x"20",x"C3", -- 0xB998
    x"00",x"00",x"DD",x"CF",x"97",x"F2",x"DC",x"20", -- 0xB9A0
    x"C3",x"00",x"00",x"DD",x"D8",x"97",x"F5",x"DC", -- 0xB9A8
    x"20",x"C3",x"00",x"00",x"DD",x"E1",x"97",x"F8", -- 0xB9B0
    x"DC",x"20",x"C3",x"00",x"00",x"DD",x"EA",x"97", -- 0xB9B8
    x"FB",x"B6",x"0A",x"00",x"BB",x"0A",x"00",x"F6", -- 0xB9C0
    x"0A",x"00",x"FB",x"0A",x"00",x"FD",x"FF",x"7A", -- 0xB9C8
    x"0A",x"B2",x"26",x"C9",x"0A",x"B3",x"26",x"B3", -- 0xB9D0
    x"0A",x"B4",x"26",x"AB",x"A6",x"28",x"97",x"B4", -- 0xB9D8
    x"37",x"06",x"97",x"B7",x"4C",x"27",x"0E",x"D7", -- 0xB9E0
    x"CD",x"37",x"06",x"97",x"D6",x"D7",x"DF",x"37", -- 0xB9E8
    x"02",x"97",x"E8",x"20",x"92",x"10",x"AE",x"A4", -- 0xB9F0
    x"26",x"03",x"7E",x"CE",x"B3",x"EC",x"23",x"97", -- 0xB9F8
    x"F1",x"D7",x"F4",x"EC",x"25",x"97",x"F7",x"D7", -- 0xBA00
    x"FA",x"A6",x"29",x"97",x"C7",x"EE",x"2A",x"20", -- 0xBA08
    x"CB",x"34",x"76",x"BD",x"DB",x"25",x"35",x"76", -- 0xBA10
    x"0F",x"53",x"0D",x"5A",x"27",x"1F",x"39",x"0C", -- 0xBA18
    x"5A",x"0F",x"5C",x"0C",x"53",x"32",x"64",x"DC", -- 0xBA20
    x"60",x"34",x"06",x"BD",x"D4",x"D8",x"AE",x"E4", -- 0xBA28
    x"BD",x"C9",x"34",x"0D",x"5A",x"27",x"03",x"BD", -- 0xBA30
    x"D8",x"69",x"7E",x"DD",x"A4",x"CE",x"00",x"0D", -- 0xBA38
    x"10",x"8E",x"00",x"46",x"8E",x"04",x"20",x"D6", -- 0xBA40
    x"69",x"34",x"04",x"CC",x"43",x"74",x"D3",x"A9", -- 0xBA48
    x"ED",x"81",x"CC",x"60",x"59",x"ED",x"81",x"CC", -- 0xBA50
    x"37",x"55",x"AB",x"A0",x"ED",x"81",x"C6",x"6B", -- 0xBA58
    x"A6",x"C1",x"2A",x"03",x"C6",x"6D",x"40",x"E7", -- 0xBA60
    x"80",x"8B",x"90",x"19",x"89",x"40",x"19",x"8A", -- 0xBA68
    x"40",x"A7",x"80",x"6A",x"E4",x"26",x"DB",x"20", -- 0xBA70
    x"C1",x"1A",x"26",x"EA",x"29",x"3B",x"2B",x"AF", -- 0xBA78
    x"2E",x"48",x"31",x"08",x"33",x"F3",x"37",x"0A", -- 0xBA80
    x"3A",x"50",x"3D",x"C8",x"41",x"74",x"45",x"58", -- 0xBA88
    x"49",x"78",x"00",x"4E",x"20",x"08",x"21",x"EF", -- 0xBA90
    x"23",x"F4",x"26",x"18",x"28",x"5C",x"2A",x"C2", -- 0xBA98
    x"2D",x"4D",x"2F",x"FF",x"32",x"D9",x"35",x"DF", -- 0xBAA0
    x"39",x"14",x"3C",x"78",x"00",x"40",x"A5",x"4A", -- 0xBAA8
    x"85",x"42",x"00",x"01",x"02",x"03",x"04",x"00", -- 0xBAB0
    x"02",x"01",x"03",x"04",x"02",x"00",x"01",x"03", -- 0xBAB8
    x"04",x"00",x"02",x"03",x"01",x"04",x"02",x"00", -- 0xBAC0
    x"03",x"01",x"04",x"02",x"03",x"00",x"01",x"04", -- 0xBAC8
    x"00",x"02",x"03",x"04",x"01",x"02",x"00",x"03", -- 0xBAD0
    x"04",x"01",x"02",x"03",x"00",x"04",x"01",x"02", -- 0xBAD8
    x"03",x"04",x"00",x"01",x"34",x"40",x"8D",x"3D", -- 0xBAE0
    x"DE",x"4F",x"EF",x"9F",x"00",x"51",x"DF",x"51", -- 0xBAE8
    x"8E",x"00",x"43",x"C6",x"03",x"BD",x"D4",x"B1", -- 0xBAF0
    x"96",x"18",x"10",x"8E",x"DA",x"B2",x"31",x"A6", -- 0xBAF8
    x"86",x"05",x"97",x"AC",x"A6",x"80",x"E6",x"A0", -- 0xBB00
    x"A7",x"C5",x"0A",x"AC",x"26",x"F6",x"33",x"45", -- 0xBB08
    x"C6",x"04",x"BD",x"D4",x"B1",x"9E",x"7A",x"CC", -- 0xBB10
    x"FF",x"0C",x"A7",x"80",x"9F",x"4F",x"3A",x"9F", -- 0xBB18
    x"4D",x"9F",x"7A",x"35",x"C0",x"9E",x"8A",x"CE", -- 0xBB20
    x"08",x"02",x"C6",x"05",x"EF",x"81",x"33",x"C8", -- 0xBB28
    x"42",x"5A",x"26",x"F8",x"0D",x"53",x"10",x"26", -- 0xBB30
    x"01",x"4E",x"10",x"9E",x"7A",x"10",x"9C",x"78", -- 0xBB38
    x"10",x"22",x"F3",x"6F",x"30",x"A8",x"1F",x"9C", -- 0xBB40
    x"5E",x"23",x"27",x"0D",x"59",x"26",x"23",x"8E", -- 0xBB48
    x"CD",x"40",x"CE",x"04",x"2E",x"BD",x"D3",x"08", -- 0xBB50
    x"33",x"41",x"DF",x"88",x"86",x"59",x"0D",x"57", -- 0xBB58
    x"26",x"03",x"BD",x"CC",x"09",x"B7",x"04",x"37", -- 0xBB60
    x"9E",x"60",x"81",x"59",x"10",x"26",x"F6",x"C3", -- 0xBB68
    x"0C",x"59",x"30",x"A9",x"00",x"A0",x"9C",x"60", -- 0xBB70
    x"10",x"24",x"F6",x"9D",x"CC",x"FF",x"05",x"34", -- 0xBB78
    x"06",x"9E",x"8A",x"A6",x"91",x"A1",x"E4",x"24", -- 0xBB80
    x"02",x"A7",x"E4",x"5A",x"26",x"F5",x"35",x"06", -- 0xBB88
    x"81",x"FF",x"10",x"27",x"00",x"EF",x"A7",x"A0", -- 0xBB90
    x"34",x"06",x"C6",x"05",x"E0",x"61",x"58",x"D7", -- 0xBB98
    x"10",x"9E",x"8A",x"3A",x"EE",x"84",x"EC",x"C4", -- 0xBBA0
    x"81",x"FF",x"27",x"0C",x"A0",x"E4",x"A7",x"C4", -- 0xBBA8
    x"26",x"04",x"33",x"42",x"EF",x"84",x"C1",x"70", -- 0xBBB0
    x"27",x"77",x"34",x"04",x"C4",x"70",x"C1",x"60", -- 0xBBB8
    x"35",x"04",x"27",x"67",x"D7",x"6B",x"C4",x"8F", -- 0xBBC0
    x"26",x"02",x"CA",x"10",x"2A",x"03",x"C8",x"7F", -- 0xBBC8
    x"5C",x"CB",x"0E",x"8E",x"00",x"0D",x"96",x"10", -- 0xBBD0
    x"EB",x"86",x"8C",x"C0",x"0E",x"CB",x"07",x"2B", -- 0xBBD8
    x"FC",x"C1",x"2A",x"24",x"F6",x"8E",x"DC",x"5B", -- 0xBBE0
    x"3A",x"34",x"10",x"C0",x"07",x"2A",x"FC",x"8E", -- 0xBBE8
    x"DC",x"5B",x"E6",x"85",x"34",x"04",x"D6",x"16", -- 0xBBF0
    x"27",x"06",x"96",x"10",x"47",x"C6",x"07",x"3D", -- 0xBBF8
    x"EB",x"E0",x"8E",x"00",x"20",x"3A",x"86",x"70", -- 0xBC00
    x"94",x"6B",x"27",x"0A",x"BD",x"CE",x"7C",x"CE", -- 0xBC08
    x"DC",x"4E",x"E6",x"C6",x"E7",x"84",x"96",x"14", -- 0xBC10
    x"AB",x"84",x"35",x"10",x"AB",x"84",x"8C",x"80", -- 0xBC18
    x"18",x"8B",x"0C",x"2F",x"FC",x"81",x"48",x"24", -- 0xBC20
    x"F6",x"20",x"07",x"1F",x"98",x"84",x"0F",x"43", -- 0xBC28
    x"21",x"4F",x"48",x"8B",x"20",x"D6",x"10",x"57", -- 0xBC30
    x"DB",x"18",x"8E",x"DA",x"B2",x"E6",x"85",x"A7", -- 0xBC38
    x"A5",x"35",x"06",x"5A",x"10",x"26",x"FF",x"50", -- 0xBC40
    x"96",x"69",x"31",x"A6",x"7E",x"DB",x"3D",x"00", -- 0xBC48
    x"01",x"02",x"FF",x"FE",x"01",x"03",x"05",x"00", -- 0xBC50
    x"02",x"04",x"06",x"F5",x"F7",x"F9",x"FA",x"FC", -- 0xBC58
    x"FE",x"00",x"01",x"03",x"05",x"06",x"08",x"0A", -- 0xBC60
    x"0C",x"0D",x"0F",x"11",x"12",x"14",x"16",x"18", -- 0xBC68
    x"19",x"1B",x"1D",x"1E",x"20",x"22",x"24",x"25", -- 0xBC70
    x"27",x"29",x"2A",x"2C",x"2E",x"30",x"31",x"33", -- 0xBC78
    x"35",x"36",x"38",x"3A",x"3C",x"10",x"9F",x"7A", -- 0xBC80
    x"86",x"06",x"97",x"AC",x"0F",x"10",x"8E",x"08", -- 0xBC88
    x"00",x"DE",x"8A",x"CC",x"FF",x"60",x"ED",x"81", -- 0xBC90
    x"0A",x"AC",x"27",x"0F",x"AF",x"C1",x"C6",x"40", -- 0xBC98
    x"A7",x"80",x"5A",x"26",x"FB",x"20",x"EC",x"A6", -- 0xBCA0
    x"80",x"A7",x"C0",x"39",x"9E",x"5E",x"1F",x"13", -- 0xBCA8
    x"8C",x"8D",x"F4",x"8D",x"F2",x"2A",x"17",x"84", -- 0xBCB0
    x"7F",x"10",x"27",x"00",x"BA",x"81",x"60",x"26", -- 0xBCB8
    x"0D",x"33",x"5F",x"6D",x"1F",x"2A",x"EC",x"69", -- 0xBCC0
    x"84",x"43",x"66",x"84",x"20",x"E5",x"81",x"6F", -- 0xBCC8
    x"27",x"10",x"81",x"4D",x"27",x"14",x"81",x"50", -- 0xBCD0
    x"27",x"D7",x"81",x"60",x"26",x"D5",x"33",x"5F", -- 0xBCD8
    x"20",x"D1",x"A6",x"84",x"2B",x"CD",x"8D",x"BF", -- 0xBCE0
    x"20",x"F8",x"A6",x"84",x"2B",x"C5",x"8D",x"B7", -- 0xBCE8
    x"81",x"60",x"27",x"BF",x"33",x"5F",x"20",x"F2", -- 0xBCF0
    x"8D",x"0E",x"E6",x"C2",x"2A",x"FA",x"0D",x"14", -- 0xBCF8
    x"27",x"49",x"8D",x"49",x"27",x"F8",x"D7",x"18", -- 0xBD00
    x"7E",x"DF",x"7C",x"0D",x"14",x"26",x"31",x"0C", -- 0xBD08
    x"14",x"CE",x"CD",x"40",x"8D",x"E4",x"D6",x"14", -- 0xBD10
    x"27",x"26",x"9E",x"5E",x"9F",x"04",x"20",x"1D", -- 0xBD18
    x"0D",x"14",x"2B",x"1C",x"39",x"0D",x"14",x"26", -- 0xBD20
    x"17",x"0A",x"14",x"20",x"04",x"0D",x"14",x"26", -- 0xBD28
    x"1A",x"BD",x"C9",x"0D",x"8E",x"10",x"64",x"9F", -- 0xBD30
    x"02",x"9F",x"12",x"E7",x"84",x"86",x"08",x"8C", -- 0xBD38
    x"DC",x"8A",x"B7",x"FF",x"22",x"D7",x"14",x"C6", -- 0xBD40
    x"0D",x"8D",x"BD",x"5F",x"39",x"BD",x"CC",x"5B", -- 0xBD48
    x"27",x"F9",x"5D",x"2B",x"07",x"C1",x"60",x"25", -- 0xBD50
    x"02",x"C0",x"40",x"39",x"58",x"27",x"C6",x"2A", -- 0xBD58
    x"AA",x"1A",x"FF",x"8D",x"E2",x"9F",x"6D",x"9E", -- 0xBD60
    x"5E",x"CE",x"10",x"64",x"11",x"93",x"02",x"24", -- 0xBD68
    x"0D",x"DF",x"5E",x"DE",x"02",x"33",x"41",x"9E", -- 0xBD70
    x"74",x"30",x"01",x"BD",x"D2",x"AC",x"BD",x"C9", -- 0xBD78
    x"2D",x"0D",x"70",x"27",x"1F",x"0F",x"70",x"FF", -- 0xBD80
    x"00",x"78",x"12",x"10",x"CE",x"00",x"FA",x"BD", -- 0xBD88
    x"CE",x"B7",x"BD",x"C9",x"08",x"9E",x"5E",x"0D", -- 0xBD90
    x"70",x"26",x"C6",x"8E",x"DD",x"8A",x"9F",x"72", -- 0xBD98
    x"C6",x"55",x"D7",x"71",x"0F",x"58",x"7E",x"CB", -- 0xBDA0
    x"E9",x"20",x"95",x"9E",x"8A",x"C6",x"19",x"BD", -- 0xBDA8
    x"C9",x"F6",x"0A",x"16",x"CC",x"08",x"02",x"97", -- 0xBDB0
    x"06",x"97",x"0A",x"4C",x"97",x"08",x"97",x"0C", -- 0xBDB8
    x"10",x"8E",x"FF",x"20",x"E7",x"A4",x"9E",x"6D", -- 0xBDC0
    x"9F",x"88",x"0C",x"70",x"7C",x"FF",x"C7",x"1C", -- 0xBDC8
    x"EF",x"0D",x"14",x"2F",x"02",x"8D",x"06",x"8D", -- 0xBDD0
    x"60",x"8D",x"4B",x"20",x"F4",x"0D",x"01",x"26", -- 0xBDD8
    x"44",x"9E",x"04",x"9C",x"74",x"22",x"C2",x"E6", -- 0xBDE0
    x"80",x"9F",x"04",x"C4",x"7F",x"27",x"BA",x"C1", -- 0xBDE8
    x"6F",x"26",x"0A",x"6D",x"1F",x"2A",x"06",x"C6", -- 0xBDF0
    x"60",x"8D",x"30",x"C6",x"6F",x"8D",x"2C",x"6D", -- 0xBDF8
    x"9F",x"00",x"04",x"2A",x"20",x"C6",x"0D",x"8D", -- 0xBE00
    x"22",x"8C",x"8D",x"2D",x"8D",x"18",x"D6",x"18", -- 0xBE08
    x"27",x"0A",x"0D",x"00",x"27",x"F6",x"E1",x"9F", -- 0xBE10
    x"00",x"06",x"26",x"EE",x"8D",x"1B",x"8D",x"06", -- 0xBE18
    x"13",x"0D",x"00",x"26",x"F7",x"39",x"BD",x"DD", -- 0xBE20
    x"4D",x"27",x"FA",x"C1",x"60",x"25",x"02",x"C0", -- 0xBE28
    x"40",x"0C",x"09",x"E7",x"9F",x"00",x"08",x"0C", -- 0xBE30
    x"01",x"D6",x"00",x"27",x"E8",x"E6",x"9F",x"00", -- 0xBE38
    x"06",x"0C",x"07",x"0A",x"00",x"C1",x"12",x"10", -- 0xBE40
    x"27",x"FE",x"E2",x"C1",x"14",x"10",x"27",x"FE", -- 0xBE48
    x"CF",x"BD",x"DF",x"7C",x"0D",x"14",x"27",x"CD", -- 0xBE50
    x"2A",x"1B",x"9E",x"02",x"9C",x"74",x"10",x"24", -- 0xBE58
    x"FE",x"DE",x"C1",x"0D",x"26",x"28",x"0F",x"15", -- 0xBE60
    x"CC",x"80",x"E0",x"A1",x"84",x"26",x"02",x"E7", -- 0xBE68
    x"80",x"9F",x"12",x"20",x"34",x"C1",x"13",x"26", -- 0xBE70
    x"14",x"BD",x"DD",x"4D",x"0D",x"14",x"2F",x"0D", -- 0xBE78
    x"DC",x"06",x"DB",x"00",x"5A",x"1F",x"01",x"E6", -- 0xBE80
    x"84",x"C1",x"11",x"26",x"EC",x"39",x"C1",x"40", -- 0xBE88
    x"25",x"FB",x"C1",x"6F",x"26",x"0E",x"0A",x"15", -- 0xBE90
    x"A6",x"1F",x"81",x"E0",x"26",x"06",x"30",x"1F", -- 0xBE98
    x"86",x"80",x"A7",x"84",x"EA",x"84",x"E7",x"80", -- 0xBEA0
    x"4F",x"A7",x"84",x"9F",x"02",x"1F",x"10",x"93", -- 0xBEA8
    x"12",x"C1",x"20",x"26",x"D8",x"E6",x"82",x"9F", -- 0xBEB0
    x"12",x"0D",x"15",x"27",x"E3",x"86",x"EF",x"A7", -- 0xBEB8
    x"80",x"6F",x"84",x"20",x"DF",x"E6",x"22",x"54", -- 0xBEC0
    x"DC",x"0E",x"2B",x"09",x"26",x"0B",x"25",x"23", -- 0xBEC8
    x"CC",x"08",x"27",x"20",x"1C",x"24",x"1C",x"20", -- 0xBED0
    x"17",x"5A",x"26",x"15",x"66",x"9F",x"00",x"0A", -- 0xBED8
    x"C6",x"1A",x"4A",x"26",x"0C",x"9E",x"0A",x"68", -- 0xBEE0
    x"84",x"5F",x"66",x"84",x"0C",x"0B",x"0C",x"00", -- 0xBEE8
    x"43",x"DD",x"0E",x"DC",x"10",x"27",x"14",x"5A", -- 0xBEF0
    x"26",x"1F",x"53",x"66",x"9F",x"00",x"0C",x"59", -- 0xBEF8
    x"59",x"C4",x"02",x"E7",x"A4",x"5F",x"4A",x"27", -- 0xBF00
    x"10",x"20",x"0C",x"0D",x"01",x"27",x"0C",x"0C", -- 0xBF08
    x"0D",x"0A",x"01",x"86",x"0B",x"6F",x"A4",x"C6", -- 0xBF10
    x"1A",x"DD",x"10",x"B6",x"FF",x"00",x"97",x"6A", -- 0xBF18
    x"3B",x"BD",x"CE",x"B7",x"DD",x"AA",x"5F",x"DD", -- 0xBF20
    x"70",x"DD",x"A8",x"DD",x"8A",x"86",x"7E",x"8E", -- 0xBF28
    x"DE",x"C5",x"CE",x"01",x"0F",x"36",x"12",x"8E", -- 0xBF30
    x"D4",x"7D",x"36",x"12",x"8D",x"33",x"0C",x"88", -- 0xBF38
    x"BD",x"DD",x"3D",x"35",x"40",x"8C",x"8D",x"34", -- 0xBF40
    x"E6",x"C0",x"2A",x"FA",x"9E",x"AD",x"A6",x"80", -- 0xBF48
    x"8A",x"40",x"A7",x"89",x"FD",x"FF",x"8C",x"08", -- 0xBF50
    x"00",x"26",x"F3",x"BD",x"CC",x"09",x"80",x"1D", -- 0xBF58
    x"97",x"B9",x"8D",x"0D",x"8E",x"C0",x"90",x"CE", -- 0xBF60
    x"C8",x"62",x"9F",x"5E",x"0C",x"70",x"7E",x"DD", -- 0xBF68
    x"77",x"8E",x"06",x"00",x"9F",x"88",x"9F",x"6D", -- 0xBF70
    x"9F",x"AD",x"20",x"78",x"8D",x"1B",x"C1",x"20", -- 0xBF78
    x"25",x"45",x"C1",x"60",x"25",x"02",x"C0",x"20", -- 0xBF80
    x"C4",x"BF",x"E7",x"80",x"CA",x"40",x"0F",x"17", -- 0xBF88
    x"0A",x"17",x"9F",x"88",x"8C",x"08",x"00",x"24", -- 0xBF90
    x"4A",x"9E",x"88",x"A6",x"84",x"88",x"40",x"A7", -- 0xBF98
    x"84",x"39",x"1E",x"10",x"C4",x"F8",x"1E",x"10", -- 0xBFA0
    x"30",x"08",x"20",x"E2",x"0C",x"16",x"27",x"E9", -- 0xBFA8
    x"0C",x"17",x"96",x"89",x"84",x"1F",x"9A",x"17", -- 0xBFB0
    x"27",x"DF",x"30",x"88",x"21",x"9C",x"AD",x"23", -- 0xBFB8
    x"D8",x"86",x"20",x"A7",x"82",x"20",x"CB",x"C1", -- 0xBFC0
    x"09",x"27",x"D7",x"C1",x"0A",x"27",x"DD",x"C1", -- 0xBFC8
    x"08",x"27",x"EA",x"C1",x"0D",x"26",x"C2",x"1E", -- 0xBFD0
    x"10",x"C4",x"E0",x"1E",x"10",x"0F",x"16",x"0A", -- 0xBFD8
    x"16",x"20",x"CD",x"30",x"88",x"E0",x"9F",x"88", -- 0xBFE0
    x"9E",x"AD",x"A6",x"88",x"20",x"A7",x"80",x"8C", -- 0xBFE8
    x"07",x"E0",x"25",x"F6",x"86",x"20",x"A7",x"80", -- 0xBFF0
    x"8C",x"08",x"00",x"25",x"F9",x"20",x"9A",x"FF", -- 0xBFF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC000
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC008
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC010
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC018
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC020
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC028
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC030
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC038
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC040
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC048
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC050
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC060
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC068
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC070
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC078
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC080
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC088
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC090
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC098
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC0F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC100
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC108
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC110
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC118
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC120
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC128
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC130
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC138
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC140
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC148
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC150
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC158
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC160
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC168
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC170
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC178
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC180
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC188
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC190
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC198
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC1F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC200
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC208
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC210
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC218
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC220
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC228
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC230
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC238
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC240
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC248
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC250
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC258
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC260
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC268
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC270
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC278
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC280
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC288
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC290
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC298
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC2F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC300
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC308
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC310
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC318
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC320
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC328
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC330
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC338
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC340
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC348
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC350
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC358
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC360
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC368
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC370
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC378
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC380
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC388
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC390
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC398
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC3F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC400
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC408
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC410
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC418
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC420
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC428
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC430
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC438
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC440
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC448
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC450
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC458
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC460
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC468
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC470
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC478
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC480
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC488
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC490
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC498
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC4F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC500
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC508
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC510
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC518
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC520
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC528
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC530
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC538
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC540
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC548
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC550
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC558
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC560
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC568
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC570
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC578
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC580
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC588
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC590
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC598
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC5F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC600
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC608
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC610
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC618
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC620
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC628
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC630
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC638
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC640
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC648
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC650
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC658
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC660
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC668
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC670
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC678
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC680
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC688
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC690
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC698
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC6F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC700
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC708
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC710
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC718
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC720
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC728
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC730
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC738
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC740
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC748
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC750
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC758
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC760
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC768
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC770
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC778
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC780
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC788
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC790
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC798
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC7F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC800
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC808
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC810
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC818
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC820
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC828
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC830
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC838
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC840
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC848
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC850
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC858
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC860
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC868
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC870
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC878
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC880
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC888
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC890
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC898
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC8F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC900
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC908
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC910
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC918
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC920
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC928
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC930
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC938
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC940
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC948
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC950
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC958
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC960
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC968
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC970
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC978
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC980
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC988
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC990
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC998
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xC9F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCA98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCAF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCB98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCBF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCC98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCCF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCD98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCDF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCE98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCEA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCEA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCEB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCEB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCEC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCEC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCED0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCEE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCEE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCEF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCEF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCF98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xCFF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD000
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD008
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD010
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD018
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD020
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD028
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD030
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD038
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD040
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD048
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD050
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD060
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD068
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD070
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD078
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD080
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD088
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD090
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD098
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD0F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD100
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD108
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD110
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD118
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD120
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD128
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD130
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD138
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD140
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD148
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD150
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD158
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD160
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD168
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD170
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD178
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD180
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD188
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD190
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD198
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD1F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD200
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD208
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD210
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD218
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD220
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD228
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD230
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD238
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD240
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD248
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD250
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD258
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD260
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD268
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD270
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD278
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD280
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD288
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD290
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD298
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD2F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD300
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD308
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD310
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD318
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD320
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD328
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD330
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD338
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD340
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD348
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD350
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD358
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD360
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD368
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD370
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD378
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD380
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD388
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD390
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD398
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD3F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD400
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD408
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD410
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD418
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD420
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD428
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD430
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD438
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD440
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD448
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD450
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD458
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD460
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD468
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD470
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD478
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD480
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD488
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD490
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD498
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD4F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD500
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD508
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD510
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD518
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD520
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD528
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD530
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD538
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD540
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD548
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD550
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD558
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD560
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD568
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD570
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD578
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD580
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD588
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD590
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD598
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD5F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD600
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD608
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD610
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD618
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD620
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD628
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD630
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD638
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD640
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD648
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD650
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD658
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD660
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD668
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD670
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD678
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD680
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD688
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD690
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD698
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD6F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD700
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD708
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD710
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD718
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD720
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD728
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD730
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD738
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD740
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD748
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD750
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD758
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD760
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD768
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD770
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD778
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD780
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD788
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD790
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD798
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD7F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD800
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD808
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD810
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD818
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD820
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD828
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD830
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD838
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD840
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD848
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD850
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD858
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD860
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD868
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD870
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD878
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD880
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD888
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD890
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD898
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD8F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD900
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD908
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD910
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD918
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD920
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD928
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD930
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD938
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD940
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD948
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD950
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD958
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD960
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD968
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD970
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD978
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD980
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD988
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD990
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD998
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xD9F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDA98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDAF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDB98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDBF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDC98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDCF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDD98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDDF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDE98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDEA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDEA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDEB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDEB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDEC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDEC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDED0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDEE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDEE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDEF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDEF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDF98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xDFF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE000
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE008
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE010
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE018
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE020
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE028
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE030
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE038
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE040
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE048
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE050
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE060
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE068
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE070
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE078
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE080
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE088
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE090
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE098
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE0F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE100
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE108
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE110
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE118
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE120
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE128
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE130
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE138
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE140
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE148
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE150
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE158
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE160
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE168
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE170
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE178
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE180
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE188
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE190
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE198
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE1F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE200
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE208
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE210
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE218
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE220
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE228
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE230
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE238
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE240
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE248
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE250
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE258
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE260
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE268
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE270
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE278
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE280
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE288
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE290
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE298
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE2F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE300
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE308
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE310
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE318
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE320
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE328
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE330
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE338
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE340
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE348
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE350
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE358
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE360
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE368
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE370
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE378
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE380
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE388
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE390
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE398
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE3F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE400
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE408
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE410
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE418
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE420
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE428
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE430
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE438
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE440
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE448
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE450
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE458
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE460
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE468
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE470
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE478
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE480
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE488
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE490
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE498
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE4F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE500
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE508
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE510
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE518
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE520
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE528
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE530
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE538
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE540
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE548
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE550
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE558
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE560
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE568
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE570
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE578
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE580
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE588
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE590
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE598
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE5F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE600
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE608
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE610
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE618
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE620
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE628
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE630
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE638
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE640
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE648
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE650
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE658
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE660
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE668
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE670
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE678
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE680
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE688
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE690
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE698
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE6F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE700
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE708
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE710
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE718
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE720
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE728
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE730
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE738
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE740
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE748
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE750
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE758
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE760
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE768
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE770
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE778
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE780
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE788
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE790
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE798
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE7F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE800
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE808
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE810
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE818
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE820
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE828
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE830
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE838
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE840
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE848
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE850
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE858
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE860
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE868
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE870
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE878
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE880
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE888
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE890
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE898
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE8F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE900
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE908
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE910
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE918
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE920
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE928
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE930
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE938
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE940
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE948
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE950
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE958
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE960
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE968
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE970
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE978
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE980
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE988
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE990
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE998
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xE9F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEA98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEAF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEB98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEBF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEC98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xECF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xED98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEDF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEE98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEEA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEEA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEEB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEEB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEEC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEEC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEED0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEEE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEEE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEEF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEEF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEF98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xEFF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF000
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF008
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF010
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF018
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF020
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF028
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF030
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF038
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF040
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF048
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF050
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF060
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF068
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF070
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF078
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF080
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF088
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF090
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF098
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF0F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF100
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF108
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF110
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF118
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF120
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF128
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF130
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF138
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF140
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF148
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF150
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF158
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF160
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF168
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF170
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF178
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF180
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF188
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF190
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF198
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF1F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF200
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF208
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF210
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF218
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF220
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF228
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF230
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF238
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF240
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF248
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF250
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF258
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF260
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF268
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF270
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF278
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF280
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF288
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF290
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF298
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF2F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF300
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF308
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF310
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF318
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF320
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF328
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF330
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF338
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF340
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF348
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF350
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF358
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF360
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF368
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF370
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF378
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF380
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF388
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF390
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF398
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF3F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF400
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF408
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF410
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF418
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF420
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF428
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF430
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF438
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF440
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF448
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF450
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF458
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF460
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF468
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF470
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF478
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF480
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF488
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF490
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF498
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF4F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF500
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF508
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF510
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF518
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF520
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF528
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF530
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF538
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF540
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF548
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF550
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF558
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF560
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF568
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF570
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF578
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF580
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF588
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF590
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF598
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF5F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF600
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF608
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF610
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF618
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF620
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF628
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF630
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF638
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF640
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF648
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF650
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF658
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF660
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF668
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF670
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF678
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF680
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF688
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF690
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF698
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF6F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF700
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF708
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF710
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF718
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF720
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF728
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF730
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF738
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF740
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF748
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF750
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF758
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF760
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF768
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF770
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF778
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF780
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF788
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF790
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF798
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF7F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF800
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF808
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF810
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF818
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF820
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF828
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF830
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF838
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF840
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF848
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF850
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF858
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF860
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF868
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF870
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF878
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF880
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF888
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF890
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF898
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF8F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF900
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF908
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF910
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF918
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF920
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF928
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF930
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF938
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF940
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF948
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF950
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF958
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF960
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF968
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF970
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF978
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF980
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF988
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF990
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF998
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xF9F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFA98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFAF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFB98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFBF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFC98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFCF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFD98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFDF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFE98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFEA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFEA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFEB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFEB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFEC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFEC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFED0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFEE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFEE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFEF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFEF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFF98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0xFFF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0xFFF8
  );

begin
dp_rom_p1: process(ADDR)
  begin
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;

  dp_rom_p2: process(CLK)
  begin
    if CLK'event and CLK='1' then
        if WR = '1' then
            ROM(to_integer(unsigned(WR_ADDR))) <= WR_DATA;
        end if;
    end if;
  end process;
  
end RTL;
